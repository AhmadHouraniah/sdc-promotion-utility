// Large Scale IP - Rewritten for clean testing// Large scale performance test IP

// This IP represents a high-performance data processing unit with wide buses// Testing with thousands of signals and deep hierarchy

module large_scale_ip (module large_scale_ip (

    // Clock and reset    // Clock and reset

    input wire sys_clk,    input clk_main_200mhz,

    input wire aux_clk,    input clk_aux_100mhz,

    input wire reset_n,    input clk_slow_25mhz,

        input reset_n,

    // Wide data buses - representing large-scale design    

    input wire [511:0] data_in_wide,    input [31:0] \input_data_bus_0000_wide_signal ,

    output wire [511:0] data_out_wide,    input [31:0] \input_data_bus_0001_wide_signal ,

        input [31:0] \input_data_bus_0002_wide_signal ,

    // Control and address buses    input [31:0] \input_data_bus_0003_wide_signal ,

    input wire [127:0] addr_bus,    input [31:0] \input_data_bus_0004_wide_signal ,

    input wire [31:0] control_bus,    input [31:0] \input_data_bus_0005_wide_signal ,

    output wire [31:0] status_bus,    input [31:0] \input_data_bus_0006_wide_signal ,

        input [31:0] \input_data_bus_0007_wide_signal ,

    // Multiple processing channels    input [31:0] \input_data_bus_0008_wide_signal ,

    input wire [63:0] channel_0_data,    input [31:0] \input_data_bus_0009_wide_signal ,

    input wire [63:0] channel_1_data,    input [31:0] \input_data_bus_0010_wide_signal ,

    input wire [63:0] channel_2_data,    input [31:0] \input_data_bus_0011_wide_signal ,

    input wire [63:0] channel_3_data,    input [31:0] \input_data_bus_0012_wide_signal ,

    output wire [63:0] channel_0_result,    input [31:0] \input_data_bus_0013_wide_signal ,

    output wire [63:0] channel_1_result,    input [31:0] \input_data_bus_0014_wide_signal ,

    output wire [63:0] channel_2_result,    input [31:0] \input_data_bus_0015_wide_signal ,

    output wire [63:0] channel_3_result,    input [31:0] \input_data_bus_0016_wide_signal ,

        input [31:0] \input_data_bus_0017_wide_signal ,

    // High-speed interface signals    input [31:0] \input_data_bus_0018_wide_signal ,

    input wire [15:0] cmd_interface,    input [31:0] \input_data_bus_0019_wide_signal ,

    input wire cmd_valid,    input [31:0] \input_data_bus_0020_wide_signal ,

    output wire cmd_ready,    input [31:0] \input_data_bus_0021_wide_signal ,

    output wire [15:0] response_interface,    input [31:0] \input_data_bus_0022_wide_signal ,

    output wire response_valid,    input [31:0] \input_data_bus_0023_wide_signal ,

    input wire response_ready,    input [31:0] \input_data_bus_0024_wide_signal ,

        input [31:0] \input_data_bus_0025_wide_signal ,

    // Memory interface - DDR-style signals    input [31:0] \input_data_bus_0026_wide_signal ,

    input wire [255:0] mem_read_data,    input [31:0] \input_data_bus_0027_wide_signal ,

    output wire [255:0] mem_write_data,    input [31:0] \input_data_bus_0028_wide_signal ,

    output wire [31:0] mem_addr,    input [31:0] \input_data_bus_0029_wide_signal ,

    output wire mem_read_enable,    input [31:0] \input_data_bus_0030_wide_signal ,

    output wire mem_write_enable,    input [31:0] \input_data_bus_0031_wide_signal ,

    input wire mem_ready,    input [31:0] \input_data_bus_0032_wide_signal ,

        input [31:0] \input_data_bus_0033_wide_signal ,

    // Error and debug signals    input [31:0] \input_data_bus_0034_wide_signal ,

    output wire [7:0] error_flags,    input [31:0] \input_data_bus_0035_wide_signal ,

    output wire [31:0] debug_counter,    input [31:0] \input_data_bus_0036_wide_signal ,

    input wire debug_enable,    input [31:0] \input_data_bus_0037_wide_signal ,

        input [31:0] \input_data_bus_0038_wide_signal ,

    // Performance monitoring    input [31:0] \input_data_bus_0039_wide_signal ,

    output wire [15:0] performance_counter_0,    input [31:0] \input_data_bus_0040_wide_signal ,

    output wire [15:0] performance_counter_1,    input [31:0] \input_data_bus_0041_wide_signal ,

    output wire [15:0] performance_counter_2,    input [31:0] \input_data_bus_0042_wide_signal ,

    output wire [15:0] performance_counter_3,    input [31:0] \input_data_bus_0043_wide_signal ,

    output wire [15:0] performance_counter_4,    input [31:0] \input_data_bus_0044_wide_signal ,

    output wire [15:0] performance_counter_5,    input [31:0] \input_data_bus_0045_wide_signal ,

    output wire [15:0] performance_counter_6,    input [31:0] \input_data_bus_0046_wide_signal ,

    output wire [15:0] performance_counter_7,    input [31:0] \input_data_bus_0047_wide_signal ,

    output wire busy,    input [31:0] \input_data_bus_0048_wide_signal ,

    output wire idle    input [31:0] \input_data_bus_0049_wide_signal ,

);    input [31:0] \input_data_bus_0050_wide_signal ,

    input [31:0] \input_data_bus_0051_wide_signal ,

    // Internal registers and logic    input [31:0] \input_data_bus_0052_wide_signal ,

    reg [511:0] internal_buffer_0;    input [31:0] \input_data_bus_0053_wide_signal ,

    reg [511:0] internal_buffer_1;    input [31:0] \input_data_bus_0054_wide_signal ,

    reg [127:0] addr_reg;    input [31:0] \input_data_bus_0055_wide_signal ,

    reg [31:0] control_reg;    input [31:0] \input_data_bus_0056_wide_signal ,

    reg [31:0] status_reg;    input [31:0] \input_data_bus_0057_wide_signal ,

        input [31:0] \input_data_bus_0058_wide_signal ,

    // Channel processing registers    input [31:0] \input_data_bus_0059_wide_signal ,

    reg [63:0] channel_regs [3:0];    input [31:0] \input_data_bus_0060_wide_signal ,

    reg [63:0] result_regs [3:0];    input [31:0] \input_data_bus_0061_wide_signal ,

        input [31:0] \input_data_bus_0062_wide_signal ,

    // Command processing    input [31:0] \input_data_bus_0063_wide_signal ,

    reg [15:0] cmd_reg;    input [31:0] \input_data_bus_0064_wide_signal ,

    reg cmd_valid_reg;    input [31:0] \input_data_bus_0065_wide_signal ,

    reg cmd_ready_reg;    input [31:0] \input_data_bus_0066_wide_signal ,

    reg [15:0] response_reg;    input [31:0] \input_data_bus_0067_wide_signal ,

    reg response_valid_reg;    input [31:0] \input_data_bus_0068_wide_signal ,

        input [31:0] \input_data_bus_0069_wide_signal ,

    // Memory interface registers    input [31:0] \input_data_bus_0070_wide_signal ,

    reg [255:0] mem_write_reg;    input [31:0] \input_data_bus_0071_wide_signal ,

    reg [31:0] mem_addr_reg;    input [31:0] \input_data_bus_0072_wide_signal ,

    reg mem_read_enable_reg;    input [31:0] \input_data_bus_0073_wide_signal ,

    reg mem_write_enable_reg;    input [31:0] \input_data_bus_0074_wide_signal ,

        input [31:0] \input_data_bus_0075_wide_signal ,

    // Error and debug registers    input [31:0] \input_data_bus_0076_wide_signal ,

    reg [7:0] error_reg;    input [31:0] \input_data_bus_0077_wide_signal ,

    reg [31:0] debug_counter_reg;    input [31:0] \input_data_bus_0078_wide_signal ,

        input [31:0] \input_data_bus_0079_wide_signal ,

    // Performance counters    input [31:0] \input_data_bus_0080_wide_signal ,

    reg [15:0] perf_counters [7:0];    input [31:0] \input_data_bus_0081_wide_signal ,

    reg busy_reg;    input [31:0] \input_data_bus_0082_wide_signal ,

    reg idle_reg;    input [31:0] \input_data_bus_0083_wide_signal ,

        input [31:0] \input_data_bus_0084_wide_signal ,

    // Main processing logic    input [31:0] \input_data_bus_0085_wide_signal ,

    always @(posedge sys_clk or negedge reset_n) begin    input [31:0] \input_data_bus_0086_wide_signal ,

        if (!reset_n) begin    input [31:0] \input_data_bus_0087_wide_signal ,

            // Reset all registers    input [31:0] \input_data_bus_0088_wide_signal ,

            internal_buffer_0 <= 512'h0;    input [31:0] \input_data_bus_0089_wide_signal ,

            internal_buffer_1 <= 512'h0;    input [31:0] \input_data_bus_0090_wide_signal ,

            addr_reg <= 128'h0;    input [31:0] \input_data_bus_0091_wide_signal ,

            control_reg <= 32'h0;    input [31:0] \input_data_bus_0092_wide_signal ,

            status_reg <= 32'h0;    input [31:0] \input_data_bus_0093_wide_signal ,

                input [31:0] \input_data_bus_0094_wide_signal ,

            for (integer i = 0; i < 4; i = i + 1) begin    input [31:0] \input_data_bus_0095_wide_signal ,

                channel_regs[i] <= 64'h0;    input [31:0] \input_data_bus_0096_wide_signal ,

                result_regs[i] <= 64'h0;    input [31:0] \input_data_bus_0097_wide_signal ,

            end    input [31:0] \input_data_bus_0098_wide_signal ,

                input [31:0] \input_data_bus_0099_wide_signal ,

            cmd_reg <= 16'h0;    input [31:0] \input_data_bus_0100_wide_signal ,

            cmd_valid_reg <= 1'b0;    input [31:0] \input_data_bus_0101_wide_signal ,

            cmd_ready_reg <= 1'b1;    input [31:0] \input_data_bus_0102_wide_signal ,

            response_reg <= 16'h0;    input [31:0] \input_data_bus_0103_wide_signal ,

            response_valid_reg <= 1'b0;    input [31:0] \input_data_bus_0104_wide_signal ,

                input [31:0] \input_data_bus_0105_wide_signal ,

            mem_write_reg <= 256'h0;    input [31:0] \input_data_bus_0106_wide_signal ,

            mem_addr_reg <= 32'h0;    input [31:0] \input_data_bus_0107_wide_signal ,

            mem_read_enable_reg <= 1'b0;    input [31:0] \input_data_bus_0108_wide_signal ,

            mem_write_enable_reg <= 1'b0;    input [31:0] \input_data_bus_0109_wide_signal ,

                input [31:0] \input_data_bus_0110_wide_signal ,

            error_reg <= 8'h0;    input [31:0] \input_data_bus_0111_wide_signal ,

            debug_counter_reg <= 32'h0;    input [31:0] \input_data_bus_0112_wide_signal ,

                input [31:0] \input_data_bus_0113_wide_signal ,

            for (integer i = 0; i < 8; i = i + 1) begin    input [31:0] \input_data_bus_0114_wide_signal ,

                perf_counters[i] <= 16'h0;    input [31:0] \input_data_bus_0115_wide_signal ,

            end    input [31:0] \input_data_bus_0116_wide_signal ,

                input [31:0] \input_data_bus_0117_wide_signal ,

            busy_reg <= 1'b0;    input [31:0] \input_data_bus_0118_wide_signal ,

            idle_reg <= 1'b1;    input [31:0] \input_data_bus_0119_wide_signal ,

        end else begin    input [31:0] \input_data_bus_0120_wide_signal ,

            // Data processing    input [31:0] \input_data_bus_0121_wide_signal ,

            internal_buffer_0 <= data_in_wide;    input [31:0] \input_data_bus_0122_wide_signal ,

            internal_buffer_1 <= internal_buffer_0;    input [31:0] \input_data_bus_0123_wide_signal ,

                input [31:0] \input_data_bus_0124_wide_signal ,

            // Address and control    input [31:0] \input_data_bus_0125_wide_signal ,

            addr_reg <= addr_bus;    input [31:0] \input_data_bus_0126_wide_signal ,

            control_reg <= control_bus;    input [31:0] \input_data_bus_0127_wide_signal ,

            status_reg <= {busy_reg, idle_reg, error_reg[5:0], perf_counters[0][15:8], perf_counters[1][15:8]};    input [31:0] \input_data_bus_0128_wide_signal ,

                input [31:0] \input_data_bus_0129_wide_signal ,

            // Channel processing    input [31:0] \input_data_bus_0130_wide_signal ,

            channel_regs[0] <= channel_0_data;    input [31:0] \input_data_bus_0131_wide_signal ,

            channel_regs[1] <= channel_1_data;    input [31:0] \input_data_bus_0132_wide_signal ,

            channel_regs[2] <= channel_2_data;    input [31:0] \input_data_bus_0133_wide_signal ,

            channel_regs[3] <= channel_3_data;    input [31:0] \input_data_bus_0134_wide_signal ,

                input [31:0] \input_data_bus_0135_wide_signal ,

            // Simple processing (add some delay)    input [31:0] \input_data_bus_0136_wide_signal ,

            result_regs[0] <= channel_regs[0] + 64'h1;    input [31:0] \input_data_bus_0137_wide_signal ,

            result_regs[1] <= channel_regs[1] + 64'h2;    input [31:0] \input_data_bus_0138_wide_signal ,

            result_regs[2] <= channel_regs[2] + 64'h3;    input [31:0] \input_data_bus_0139_wide_signal ,

            result_regs[3] <= channel_regs[3] + 64'h4;    input [31:0] \input_data_bus_0140_wide_signal ,

                input [31:0] \input_data_bus_0141_wide_signal ,

            // Command processing    input [31:0] \input_data_bus_0142_wide_signal ,

            if (cmd_valid && cmd_ready_reg) begin    input [31:0] \input_data_bus_0143_wide_signal ,

                cmd_reg <= cmd_interface;    input [31:0] \input_data_bus_0144_wide_signal ,

                cmd_valid_reg <= 1'b1;    input [31:0] \input_data_bus_0145_wide_signal ,

                cmd_ready_reg <= 1'b0;    input [31:0] \input_data_bus_0146_wide_signal ,

                response_reg <= cmd_interface + 16'h100; // Simple response    input [31:0] \input_data_bus_0147_wide_signal ,

                response_valid_reg <= 1'b1;    input [31:0] \input_data_bus_0148_wide_signal ,

            end    input [31:0] \input_data_bus_0149_wide_signal ,

                input [31:0] \input_data_bus_0150_wide_signal ,

            if (response_valid_reg && response_ready) begin    input [31:0] \input_data_bus_0151_wide_signal ,

                response_valid_reg <= 1'b0;    input [31:0] \input_data_bus_0152_wide_signal ,

                cmd_ready_reg <= 1'b1;    input [31:0] \input_data_bus_0153_wide_signal ,

            end    input [31:0] \input_data_bus_0154_wide_signal ,

                input [31:0] \input_data_bus_0155_wide_signal ,

            // Memory interface    input [31:0] \input_data_bus_0156_wide_signal ,

            if (control_reg[0]) begin // Read operation    input [31:0] \input_data_bus_0157_wide_signal ,

                mem_addr_reg <= addr_reg[31:0];    input [31:0] \input_data_bus_0158_wide_signal ,

                mem_read_enable_reg <= 1'b1;    input [31:0] \input_data_bus_0159_wide_signal ,

                mem_write_enable_reg <= 1'b0;    input [31:0] \input_data_bus_0160_wide_signal ,

            end else if (control_reg[1]) begin // Write operation    input [31:0] \input_data_bus_0161_wide_signal ,

                mem_addr_reg <= addr_reg[31:0];    input [31:0] \input_data_bus_0162_wide_signal ,

                mem_write_reg <= internal_buffer_1[255:0];    input [31:0] \input_data_bus_0163_wide_signal ,

                mem_write_enable_reg <= 1'b1;    input [31:0] \input_data_bus_0164_wide_signal ,

                mem_read_enable_reg <= 1'b0;    input [31:0] \input_data_bus_0165_wide_signal ,

            end else begin    input [31:0] \input_data_bus_0166_wide_signal ,

                mem_read_enable_reg <= 1'b0;    input [31:0] \input_data_bus_0167_wide_signal ,

                mem_write_enable_reg <= 1'b0;    input [31:0] \input_data_bus_0168_wide_signal ,

            end    input [31:0] \input_data_bus_0169_wide_signal ,

                input [31:0] \input_data_bus_0170_wide_signal ,

            // Debug counter    input [31:0] \input_data_bus_0171_wide_signal ,

            if (debug_enable) begin    input [31:0] \input_data_bus_0172_wide_signal ,

                debug_counter_reg <= debug_counter_reg + 32'h1;    input [31:0] \input_data_bus_0173_wide_signal ,

            end    input [31:0] \input_data_bus_0174_wide_signal ,

                input [31:0] \input_data_bus_0175_wide_signal ,

            // Performance counters    input [31:0] \input_data_bus_0176_wide_signal ,

            perf_counters[0] <= perf_counters[0] + (busy_reg ? 16'h1 : 16'h0);    input [31:0] \input_data_bus_0177_wide_signal ,

            perf_counters[1] <= perf_counters[1] + (idle_reg ? 16'h1 : 16'h0);    input [31:0] \input_data_bus_0178_wide_signal ,

            perf_counters[2] <= perf_counters[2] + (mem_read_enable_reg ? 16'h1 : 16'h0);    input [31:0] \input_data_bus_0179_wide_signal ,

            perf_counters[3] <= perf_counters[3] + (mem_write_enable_reg ? 16'h1 : 16'h0);    input [31:0] \input_data_bus_0180_wide_signal ,

            perf_counters[4] <= perf_counters[4] + (cmd_valid_reg ? 16'h1 : 16'h0);    input [31:0] \input_data_bus_0181_wide_signal ,

            perf_counters[5] <= perf_counters[5] + (response_valid_reg ? 16'h1 : 16'h0);    input [31:0] \input_data_bus_0182_wide_signal ,

            perf_counters[6] <= perf_counters[6] + (|error_reg ? 16'h1 : 16'h0);    input [31:0] \input_data_bus_0183_wide_signal ,

            perf_counters[7] <= debug_counter_reg[15:0];    input [31:0] \input_data_bus_0184_wide_signal ,

                input [31:0] \input_data_bus_0185_wide_signal ,

            // Status logic    input [31:0] \input_data_bus_0186_wide_signal ,

            busy_reg <= |control_reg[3:0] || cmd_valid_reg || mem_read_enable_reg || mem_write_enable_reg;    input [31:0] \input_data_bus_0187_wide_signal ,

            idle_reg <= !busy_reg;    input [31:0] \input_data_bus_0188_wide_signal ,

                input [31:0] \input_data_bus_0189_wide_signal ,

            // Error detection    input [31:0] \input_data_bus_0190_wide_signal ,

            if (control_reg[31]) begin // Error injection for testing    input [31:0] \input_data_bus_0191_wide_signal ,

                error_reg <= error_reg | 8'h1;    input [31:0] \input_data_bus_0192_wide_signal ,

            end    input [31:0] \input_data_bus_0193_wide_signal ,

        end    input [31:0] \input_data_bus_0194_wide_signal ,

    end    input [31:0] \input_data_bus_0195_wide_signal ,

        input [31:0] \input_data_bus_0196_wide_signal ,

    // Output assignments    input [31:0] \input_data_bus_0197_wide_signal ,

    assign data_out_wide = internal_buffer_1;    input [31:0] \input_data_bus_0198_wide_signal ,

    assign status_bus = status_reg;    input [31:0] \input_data_bus_0199_wide_signal ,

        input [31:0] \input_data_bus_0200_wide_signal ,

    assign channel_0_result = result_regs[0];    input [31:0] \input_data_bus_0201_wide_signal ,

    assign channel_1_result = result_regs[1];    input [31:0] \input_data_bus_0202_wide_signal ,

    assign channel_2_result = result_regs[2];    input [31:0] \input_data_bus_0203_wide_signal ,

    assign channel_3_result = result_regs[3];    input [31:0] \input_data_bus_0204_wide_signal ,

        input [31:0] \input_data_bus_0205_wide_signal ,

    assign cmd_ready = cmd_ready_reg;    input [31:0] \input_data_bus_0206_wide_signal ,

    assign response_interface = response_reg;    input [31:0] \input_data_bus_0207_wide_signal ,

    assign response_valid = response_valid_reg;    input [31:0] \input_data_bus_0208_wide_signal ,

        input [31:0] \input_data_bus_0209_wide_signal ,

    assign mem_write_data = mem_write_reg;    input [31:0] \input_data_bus_0210_wide_signal ,

    assign mem_addr = mem_addr_reg;    input [31:0] \input_data_bus_0211_wide_signal ,

    assign mem_read_enable = mem_read_enable_reg;    input [31:0] \input_data_bus_0212_wide_signal ,

    assign mem_write_enable = mem_write_enable_reg;    input [31:0] \input_data_bus_0213_wide_signal ,

        input [31:0] \input_data_bus_0214_wide_signal ,

    assign error_flags = error_reg;    input [31:0] \input_data_bus_0215_wide_signal ,

    assign debug_counter = debug_counter_reg;    input [31:0] \input_data_bus_0216_wide_signal ,

        input [31:0] \input_data_bus_0217_wide_signal ,

    // Performance counter outputs    input [31:0] \input_data_bus_0218_wide_signal ,

    assign performance_counter_0 = perf_counters[0];    input [31:0] \input_data_bus_0219_wide_signal ,

    assign performance_counter_1 = perf_counters[1];    input [31:0] \input_data_bus_0220_wide_signal ,

    assign performance_counter_2 = perf_counters[2];    input [31:0] \input_data_bus_0221_wide_signal ,

    assign performance_counter_3 = perf_counters[3];    input [31:0] \input_data_bus_0222_wide_signal ,

    assign performance_counter_4 = perf_counters[4];    input [31:0] \input_data_bus_0223_wide_signal ,

    assign performance_counter_5 = perf_counters[5];    input [31:0] \input_data_bus_0224_wide_signal ,

    assign performance_counter_6 = perf_counters[6];    input [31:0] \input_data_bus_0225_wide_signal ,

    assign performance_counter_7 = perf_counters[7];    input [31:0] \input_data_bus_0226_wide_signal ,

        input [31:0] \input_data_bus_0227_wide_signal ,

    assign busy = busy_reg;    input [31:0] \input_data_bus_0228_wide_signal ,

    assign idle = idle_reg;    input [31:0] \input_data_bus_0229_wide_signal ,

    input [31:0] \input_data_bus_0230_wide_signal ,

endmodule    input [31:0] \input_data_bus_0231_wide_signal ,
    input [31:0] \input_data_bus_0232_wide_signal ,
    input [31:0] \input_data_bus_0233_wide_signal ,
    input [31:0] \input_data_bus_0234_wide_signal ,
    input [31:0] \input_data_bus_0235_wide_signal ,
    input [31:0] \input_data_bus_0236_wide_signal ,
    input [31:0] \input_data_bus_0237_wide_signal ,
    input [31:0] \input_data_bus_0238_wide_signal ,
    input [31:0] \input_data_bus_0239_wide_signal ,
    input [31:0] \input_data_bus_0240_wide_signal ,
    input [31:0] \input_data_bus_0241_wide_signal ,
    input [31:0] \input_data_bus_0242_wide_signal ,
    input [31:0] \input_data_bus_0243_wide_signal ,
    input [31:0] \input_data_bus_0244_wide_signal ,
    input [31:0] \input_data_bus_0245_wide_signal ,
    input [31:0] \input_data_bus_0246_wide_signal ,
    input [31:0] \input_data_bus_0247_wide_signal ,
    input [31:0] \input_data_bus_0248_wide_signal ,
    input [31:0] \input_data_bus_0249_wide_signal ,
    input [31:0] \input_data_bus_0250_wide_signal ,
    input [31:0] \input_data_bus_0251_wide_signal ,
    input [31:0] \input_data_bus_0252_wide_signal ,
    input [31:0] \input_data_bus_0253_wide_signal ,
    input [31:0] \input_data_bus_0254_wide_signal ,
    input [31:0] \input_data_bus_0255_wide_signal ,
    input [31:0] \input_data_bus_0256_wide_signal ,
    input [31:0] \input_data_bus_0257_wide_signal ,
    input [31:0] \input_data_bus_0258_wide_signal ,
    input [31:0] \input_data_bus_0259_wide_signal ,
    input [31:0] \input_data_bus_0260_wide_signal ,
    input [31:0] \input_data_bus_0261_wide_signal ,
    input [31:0] \input_data_bus_0262_wide_signal ,
    input [31:0] \input_data_bus_0263_wide_signal ,
    input [31:0] \input_data_bus_0264_wide_signal ,
    input [31:0] \input_data_bus_0265_wide_signal ,
    input [31:0] \input_data_bus_0266_wide_signal ,
    input [31:0] \input_data_bus_0267_wide_signal ,
    input [31:0] \input_data_bus_0268_wide_signal ,
    input [31:0] \input_data_bus_0269_wide_signal ,
    input [31:0] \input_data_bus_0270_wide_signal ,
    input [31:0] \input_data_bus_0271_wide_signal ,
    input [31:0] \input_data_bus_0272_wide_signal ,
    input [31:0] \input_data_bus_0273_wide_signal ,
    input [31:0] \input_data_bus_0274_wide_signal ,
    input [31:0] \input_data_bus_0275_wide_signal ,
    input [31:0] \input_data_bus_0276_wide_signal ,
    input [31:0] \input_data_bus_0277_wide_signal ,
    input [31:0] \input_data_bus_0278_wide_signal ,
    input [31:0] \input_data_bus_0279_wide_signal ,
    input [31:0] \input_data_bus_0280_wide_signal ,
    input [31:0] \input_data_bus_0281_wide_signal ,
    input [31:0] \input_data_bus_0282_wide_signal ,
    input [31:0] \input_data_bus_0283_wide_signal ,
    input [31:0] \input_data_bus_0284_wide_signal ,
    input [31:0] \input_data_bus_0285_wide_signal ,
    input [31:0] \input_data_bus_0286_wide_signal ,
    input [31:0] \input_data_bus_0287_wide_signal ,
    input [31:0] \input_data_bus_0288_wide_signal ,
    input [31:0] \input_data_bus_0289_wide_signal ,
    input [31:0] \input_data_bus_0290_wide_signal ,
    input [31:0] \input_data_bus_0291_wide_signal ,
    input [31:0] \input_data_bus_0292_wide_signal ,
    input [31:0] \input_data_bus_0293_wide_signal ,
    input [31:0] \input_data_bus_0294_wide_signal ,
    input [31:0] \input_data_bus_0295_wide_signal ,
    input [31:0] \input_data_bus_0296_wide_signal ,
    input [31:0] \input_data_bus_0297_wide_signal ,
    input [31:0] \input_data_bus_0298_wide_signal ,
    input [31:0] \input_data_bus_0299_wide_signal ,
    input [31:0] \input_data_bus_0300_wide_signal ,
    input [31:0] \input_data_bus_0301_wide_signal ,
    input [31:0] \input_data_bus_0302_wide_signal ,
    input [31:0] \input_data_bus_0303_wide_signal ,
    input [31:0] \input_data_bus_0304_wide_signal ,
    input [31:0] \input_data_bus_0305_wide_signal ,
    input [31:0] \input_data_bus_0306_wide_signal ,
    input [31:0] \input_data_bus_0307_wide_signal ,
    input [31:0] \input_data_bus_0308_wide_signal ,
    input [31:0] \input_data_bus_0309_wide_signal ,
    input [31:0] \input_data_bus_0310_wide_signal ,
    input [31:0] \input_data_bus_0311_wide_signal ,
    input [31:0] \input_data_bus_0312_wide_signal ,
    input [31:0] \input_data_bus_0313_wide_signal ,
    input [31:0] \input_data_bus_0314_wide_signal ,
    input [31:0] \input_data_bus_0315_wide_signal ,
    input [31:0] \input_data_bus_0316_wide_signal ,
    input [31:0] \input_data_bus_0317_wide_signal ,
    input [31:0] \input_data_bus_0318_wide_signal ,
    input [31:0] \input_data_bus_0319_wide_signal ,
    input [31:0] \input_data_bus_0320_wide_signal ,
    input [31:0] \input_data_bus_0321_wide_signal ,
    input [31:0] \input_data_bus_0322_wide_signal ,
    input [31:0] \input_data_bus_0323_wide_signal ,
    input [31:0] \input_data_bus_0324_wide_signal ,
    input [31:0] \input_data_bus_0325_wide_signal ,
    input [31:0] \input_data_bus_0326_wide_signal ,
    input [31:0] \input_data_bus_0327_wide_signal ,
    input [31:0] \input_data_bus_0328_wide_signal ,
    input [31:0] \input_data_bus_0329_wide_signal ,
    input [31:0] \input_data_bus_0330_wide_signal ,
    input [31:0] \input_data_bus_0331_wide_signal ,
    input [31:0] \input_data_bus_0332_wide_signal ,
    input [31:0] \input_data_bus_0333_wide_signal ,
    input [31:0] \input_data_bus_0334_wide_signal ,
    input [31:0] \input_data_bus_0335_wide_signal ,
    input [31:0] \input_data_bus_0336_wide_signal ,
    input [31:0] \input_data_bus_0337_wide_signal ,
    input [31:0] \input_data_bus_0338_wide_signal ,
    input [31:0] \input_data_bus_0339_wide_signal ,
    input [31:0] \input_data_bus_0340_wide_signal ,
    input [31:0] \input_data_bus_0341_wide_signal ,
    input [31:0] \input_data_bus_0342_wide_signal ,
    input [31:0] \input_data_bus_0343_wide_signal ,
    input [31:0] \input_data_bus_0344_wide_signal ,
    input [31:0] \input_data_bus_0345_wide_signal ,
    input [31:0] \input_data_bus_0346_wide_signal ,
    input [31:0] \input_data_bus_0347_wide_signal ,
    input [31:0] \input_data_bus_0348_wide_signal ,
    input [31:0] \input_data_bus_0349_wide_signal ,
    input [31:0] \input_data_bus_0350_wide_signal ,
    input [31:0] \input_data_bus_0351_wide_signal ,
    input [31:0] \input_data_bus_0352_wide_signal ,
    input [31:0] \input_data_bus_0353_wide_signal ,
    input [31:0] \input_data_bus_0354_wide_signal ,
    input [31:0] \input_data_bus_0355_wide_signal ,
    input [31:0] \input_data_bus_0356_wide_signal ,
    input [31:0] \input_data_bus_0357_wide_signal ,
    input [31:0] \input_data_bus_0358_wide_signal ,
    input [31:0] \input_data_bus_0359_wide_signal ,
    input [31:0] \input_data_bus_0360_wide_signal ,
    input [31:0] \input_data_bus_0361_wide_signal ,
    input [31:0] \input_data_bus_0362_wide_signal ,
    input [31:0] \input_data_bus_0363_wide_signal ,
    input [31:0] \input_data_bus_0364_wide_signal ,
    input [31:0] \input_data_bus_0365_wide_signal ,
    input [31:0] \input_data_bus_0366_wide_signal ,
    input [31:0] \input_data_bus_0367_wide_signal ,
    input [31:0] \input_data_bus_0368_wide_signal ,
    input [31:0] \input_data_bus_0369_wide_signal ,
    input [31:0] \input_data_bus_0370_wide_signal ,
    input [31:0] \input_data_bus_0371_wide_signal ,
    input [31:0] \input_data_bus_0372_wide_signal ,
    input [31:0] \input_data_bus_0373_wide_signal ,
    input [31:0] \input_data_bus_0374_wide_signal ,
    input [31:0] \input_data_bus_0375_wide_signal ,
    input [31:0] \input_data_bus_0376_wide_signal ,
    input [31:0] \input_data_bus_0377_wide_signal ,
    input [31:0] \input_data_bus_0378_wide_signal ,
    input [31:0] \input_data_bus_0379_wide_signal ,
    input [31:0] \input_data_bus_0380_wide_signal ,
    input [31:0] \input_data_bus_0381_wide_signal ,
    input [31:0] \input_data_bus_0382_wide_signal ,
    input [31:0] \input_data_bus_0383_wide_signal ,
    input [31:0] \input_data_bus_0384_wide_signal ,
    input [31:0] \input_data_bus_0385_wide_signal ,
    input [31:0] \input_data_bus_0386_wide_signal ,
    input [31:0] \input_data_bus_0387_wide_signal ,
    input [31:0] \input_data_bus_0388_wide_signal ,
    input [31:0] \input_data_bus_0389_wide_signal ,
    input [31:0] \input_data_bus_0390_wide_signal ,
    input [31:0] \input_data_bus_0391_wide_signal ,
    input [31:0] \input_data_bus_0392_wide_signal ,
    input [31:0] \input_data_bus_0393_wide_signal ,
    input [31:0] \input_data_bus_0394_wide_signal ,
    input [31:0] \input_data_bus_0395_wide_signal ,
    input [31:0] \input_data_bus_0396_wide_signal ,
    input [31:0] \input_data_bus_0397_wide_signal ,
    input [31:0] \input_data_bus_0398_wide_signal ,
    input [31:0] \input_data_bus_0399_wide_signal ,
    input [31:0] \input_data_bus_0400_wide_signal ,
    input [31:0] \input_data_bus_0401_wide_signal ,
    input [31:0] \input_data_bus_0402_wide_signal ,
    input [31:0] \input_data_bus_0403_wide_signal ,
    input [31:0] \input_data_bus_0404_wide_signal ,
    input [31:0] \input_data_bus_0405_wide_signal ,
    input [31:0] \input_data_bus_0406_wide_signal ,
    input [31:0] \input_data_bus_0407_wide_signal ,
    input [31:0] \input_data_bus_0408_wide_signal ,
    input [31:0] \input_data_bus_0409_wide_signal ,
    input [31:0] \input_data_bus_0410_wide_signal ,
    input [31:0] \input_data_bus_0411_wide_signal ,
    input [31:0] \input_data_bus_0412_wide_signal ,
    input [31:0] \input_data_bus_0413_wide_signal ,
    input [31:0] \input_data_bus_0414_wide_signal ,
    input [31:0] \input_data_bus_0415_wide_signal ,
    input [31:0] \input_data_bus_0416_wide_signal ,
    input [31:0] \input_data_bus_0417_wide_signal ,
    input [31:0] \input_data_bus_0418_wide_signal ,
    input [31:0] \input_data_bus_0419_wide_signal ,
    input [31:0] \input_data_bus_0420_wide_signal ,
    input [31:0] \input_data_bus_0421_wide_signal ,
    input [31:0] \input_data_bus_0422_wide_signal ,
    input [31:0] \input_data_bus_0423_wide_signal ,
    input [31:0] \input_data_bus_0424_wide_signal ,
    input [31:0] \input_data_bus_0425_wide_signal ,
    input [31:0] \input_data_bus_0426_wide_signal ,
    input [31:0] \input_data_bus_0427_wide_signal ,
    input [31:0] \input_data_bus_0428_wide_signal ,
    input [31:0] \input_data_bus_0429_wide_signal ,
    input [31:0] \input_data_bus_0430_wide_signal ,
    input [31:0] \input_data_bus_0431_wide_signal ,
    input [31:0] \input_data_bus_0432_wide_signal ,
    input [31:0] \input_data_bus_0433_wide_signal ,
    input [31:0] \input_data_bus_0434_wide_signal ,
    input [31:0] \input_data_bus_0435_wide_signal ,
    input [31:0] \input_data_bus_0436_wide_signal ,
    input [31:0] \input_data_bus_0437_wide_signal ,
    input [31:0] \input_data_bus_0438_wide_signal ,
    input [31:0] \input_data_bus_0439_wide_signal ,
    input [31:0] \input_data_bus_0440_wide_signal ,
    input [31:0] \input_data_bus_0441_wide_signal ,
    input [31:0] \input_data_bus_0442_wide_signal ,
    input [31:0] \input_data_bus_0443_wide_signal ,
    input [31:0] \input_data_bus_0444_wide_signal ,
    input [31:0] \input_data_bus_0445_wide_signal ,
    input [31:0] \input_data_bus_0446_wide_signal ,
    input [31:0] \input_data_bus_0447_wide_signal ,
    input [31:0] \input_data_bus_0448_wide_signal ,
    input [31:0] \input_data_bus_0449_wide_signal ,
    input [31:0] \input_data_bus_0450_wide_signal ,
    input [31:0] \input_data_bus_0451_wide_signal ,
    input [31:0] \input_data_bus_0452_wide_signal ,
    input [31:0] \input_data_bus_0453_wide_signal ,
    input [31:0] \input_data_bus_0454_wide_signal ,
    input [31:0] \input_data_bus_0455_wide_signal ,
    input [31:0] \input_data_bus_0456_wide_signal ,
    input [31:0] \input_data_bus_0457_wide_signal ,
    input [31:0] \input_data_bus_0458_wide_signal ,
    input [31:0] \input_data_bus_0459_wide_signal ,
    input [31:0] \input_data_bus_0460_wide_signal ,
    input [31:0] \input_data_bus_0461_wide_signal ,
    input [31:0] \input_data_bus_0462_wide_signal ,
    input [31:0] \input_data_bus_0463_wide_signal ,
    input [31:0] \input_data_bus_0464_wide_signal ,
    input [31:0] \input_data_bus_0465_wide_signal ,
    input [31:0] \input_data_bus_0466_wide_signal ,
    input [31:0] \input_data_bus_0467_wide_signal ,
    input [31:0] \input_data_bus_0468_wide_signal ,
    input [31:0] \input_data_bus_0469_wide_signal ,
    input [31:0] \input_data_bus_0470_wide_signal ,
    input [31:0] \input_data_bus_0471_wide_signal ,
    input [31:0] \input_data_bus_0472_wide_signal ,
    input [31:0] \input_data_bus_0473_wide_signal ,
    input [31:0] \input_data_bus_0474_wide_signal ,
    input [31:0] \input_data_bus_0475_wide_signal ,
    input [31:0] \input_data_bus_0476_wide_signal ,
    input [31:0] \input_data_bus_0477_wide_signal ,
    input [31:0] \input_data_bus_0478_wide_signal ,
    input [31:0] \input_data_bus_0479_wide_signal ,
    input [31:0] \input_data_bus_0480_wide_signal ,
    input [31:0] \input_data_bus_0481_wide_signal ,
    input [31:0] \input_data_bus_0482_wide_signal ,
    input [31:0] \input_data_bus_0483_wide_signal ,
    input [31:0] \input_data_bus_0484_wide_signal ,
    input [31:0] \input_data_bus_0485_wide_signal ,
    input [31:0] \input_data_bus_0486_wide_signal ,
    input [31:0] \input_data_bus_0487_wide_signal ,
    input [31:0] \input_data_bus_0488_wide_signal ,
    input [31:0] \input_data_bus_0489_wide_signal ,
    input [31:0] \input_data_bus_0490_wide_signal ,
    input [31:0] \input_data_bus_0491_wide_signal ,
    input [31:0] \input_data_bus_0492_wide_signal ,
    input [31:0] \input_data_bus_0493_wide_signal ,
    input [31:0] \input_data_bus_0494_wide_signal ,
    input [31:0] \input_data_bus_0495_wide_signal ,
    input [31:0] \input_data_bus_0496_wide_signal ,
    input [31:0] \input_data_bus_0497_wide_signal ,
    input [31:0] \input_data_bus_0498_wide_signal ,
    input [31:0] \input_data_bus_0499_wide_signal ,
    input [31:0] \input_data_bus_0500_wide_signal ,
    input [31:0] \input_data_bus_0501_wide_signal ,
    input [31:0] \input_data_bus_0502_wide_signal ,
    input [31:0] \input_data_bus_0503_wide_signal ,
    input [31:0] \input_data_bus_0504_wide_signal ,
    input [31:0] \input_data_bus_0505_wide_signal ,
    input [31:0] \input_data_bus_0506_wide_signal ,
    input [31:0] \input_data_bus_0507_wide_signal ,
    input [31:0] \input_data_bus_0508_wide_signal ,
    input [31:0] \input_data_bus_0509_wide_signal ,
    input [31:0] \input_data_bus_0510_wide_signal ,
    input [31:0] \input_data_bus_0511_wide_signal ,
    input [31:0] \input_data_bus_0512_wide_signal ,
    input [31:0] \input_data_bus_0513_wide_signal ,
    input [31:0] \input_data_bus_0514_wide_signal ,
    input [31:0] \input_data_bus_0515_wide_signal ,
    input [31:0] \input_data_bus_0516_wide_signal ,
    input [31:0] \input_data_bus_0517_wide_signal ,
    input [31:0] \input_data_bus_0518_wide_signal ,
    input [31:0] \input_data_bus_0519_wide_signal ,
    input [31:0] \input_data_bus_0520_wide_signal ,
    input [31:0] \input_data_bus_0521_wide_signal ,
    input [31:0] \input_data_bus_0522_wide_signal ,
    input [31:0] \input_data_bus_0523_wide_signal ,
    input [31:0] \input_data_bus_0524_wide_signal ,
    input [31:0] \input_data_bus_0525_wide_signal ,
    input [31:0] \input_data_bus_0526_wide_signal ,
    input [31:0] \input_data_bus_0527_wide_signal ,
    input [31:0] \input_data_bus_0528_wide_signal ,
    input [31:0] \input_data_bus_0529_wide_signal ,
    input [31:0] \input_data_bus_0530_wide_signal ,
    input [31:0] \input_data_bus_0531_wide_signal ,
    input [31:0] \input_data_bus_0532_wide_signal ,
    input [31:0] \input_data_bus_0533_wide_signal ,
    input [31:0] \input_data_bus_0534_wide_signal ,
    input [31:0] \input_data_bus_0535_wide_signal ,
    input [31:0] \input_data_bus_0536_wide_signal ,
    input [31:0] \input_data_bus_0537_wide_signal ,
    input [31:0] \input_data_bus_0538_wide_signal ,
    input [31:0] \input_data_bus_0539_wide_signal ,
    input [31:0] \input_data_bus_0540_wide_signal ,
    input [31:0] \input_data_bus_0541_wide_signal ,
    input [31:0] \input_data_bus_0542_wide_signal ,
    input [31:0] \input_data_bus_0543_wide_signal ,
    input [31:0] \input_data_bus_0544_wide_signal ,
    input [31:0] \input_data_bus_0545_wide_signal ,
    input [31:0] \input_data_bus_0546_wide_signal ,
    input [31:0] \input_data_bus_0547_wide_signal ,
    input [31:0] \input_data_bus_0548_wide_signal ,
    input [31:0] \input_data_bus_0549_wide_signal ,
    input [31:0] \input_data_bus_0550_wide_signal ,
    input [31:0] \input_data_bus_0551_wide_signal ,
    input [31:0] \input_data_bus_0552_wide_signal ,
    input [31:0] \input_data_bus_0553_wide_signal ,
    input [31:0] \input_data_bus_0554_wide_signal ,
    input [31:0] \input_data_bus_0555_wide_signal ,
    input [31:0] \input_data_bus_0556_wide_signal ,
    input [31:0] \input_data_bus_0557_wide_signal ,
    input [31:0] \input_data_bus_0558_wide_signal ,
    input [31:0] \input_data_bus_0559_wide_signal ,
    input [31:0] \input_data_bus_0560_wide_signal ,
    input [31:0] \input_data_bus_0561_wide_signal ,
    input [31:0] \input_data_bus_0562_wide_signal ,
    input [31:0] \input_data_bus_0563_wide_signal ,
    input [31:0] \input_data_bus_0564_wide_signal ,
    input [31:0] \input_data_bus_0565_wide_signal ,
    input [31:0] \input_data_bus_0566_wide_signal ,
    input [31:0] \input_data_bus_0567_wide_signal ,
    input [31:0] \input_data_bus_0568_wide_signal ,
    input [31:0] \input_data_bus_0569_wide_signal ,
    input [31:0] \input_data_bus_0570_wide_signal ,
    input [31:0] \input_data_bus_0571_wide_signal ,
    input [31:0] \input_data_bus_0572_wide_signal ,
    input [31:0] \input_data_bus_0573_wide_signal ,
    input [31:0] \input_data_bus_0574_wide_signal ,
    input [31:0] \input_data_bus_0575_wide_signal ,
    input [31:0] \input_data_bus_0576_wide_signal ,
    input [31:0] \input_data_bus_0577_wide_signal ,
    input [31:0] \input_data_bus_0578_wide_signal ,
    input [31:0] \input_data_bus_0579_wide_signal ,
    input [31:0] \input_data_bus_0580_wide_signal ,
    input [31:0] \input_data_bus_0581_wide_signal ,
    input [31:0] \input_data_bus_0582_wide_signal ,
    input [31:0] \input_data_bus_0583_wide_signal ,
    input [31:0] \input_data_bus_0584_wide_signal ,
    input [31:0] \input_data_bus_0585_wide_signal ,
    input [31:0] \input_data_bus_0586_wide_signal ,
    input [31:0] \input_data_bus_0587_wide_signal ,
    input [31:0] \input_data_bus_0588_wide_signal ,
    input [31:0] \input_data_bus_0589_wide_signal ,
    input [31:0] \input_data_bus_0590_wide_signal ,
    input [31:0] \input_data_bus_0591_wide_signal ,
    input [31:0] \input_data_bus_0592_wide_signal ,
    input [31:0] \input_data_bus_0593_wide_signal ,
    input [31:0] \input_data_bus_0594_wide_signal ,
    input [31:0] \input_data_bus_0595_wide_signal ,
    input [31:0] \input_data_bus_0596_wide_signal ,
    input [31:0] \input_data_bus_0597_wide_signal ,
    input [31:0] \input_data_bus_0598_wide_signal ,
    input [31:0] \input_data_bus_0599_wide_signal ,
    input [31:0] \input_data_bus_0600_wide_signal ,
    input [31:0] \input_data_bus_0601_wide_signal ,
    input [31:0] \input_data_bus_0602_wide_signal ,
    input [31:0] \input_data_bus_0603_wide_signal ,
    input [31:0] \input_data_bus_0604_wide_signal ,
    input [31:0] \input_data_bus_0605_wide_signal ,
    input [31:0] \input_data_bus_0606_wide_signal ,
    input [31:0] \input_data_bus_0607_wide_signal ,
    input [31:0] \input_data_bus_0608_wide_signal ,
    input [31:0] \input_data_bus_0609_wide_signal ,
    input [31:0] \input_data_bus_0610_wide_signal ,
    input [31:0] \input_data_bus_0611_wide_signal ,
    input [31:0] \input_data_bus_0612_wide_signal ,
    input [31:0] \input_data_bus_0613_wide_signal ,
    input [31:0] \input_data_bus_0614_wide_signal ,
    input [31:0] \input_data_bus_0615_wide_signal ,
    input [31:0] \input_data_bus_0616_wide_signal ,
    input [31:0] \input_data_bus_0617_wide_signal ,
    input [31:0] \input_data_bus_0618_wide_signal ,
    input [31:0] \input_data_bus_0619_wide_signal ,
    input [31:0] \input_data_bus_0620_wide_signal ,
    input [31:0] \input_data_bus_0621_wide_signal ,
    input [31:0] \input_data_bus_0622_wide_signal ,
    input [31:0] \input_data_bus_0623_wide_signal ,
    input [31:0] \input_data_bus_0624_wide_signal ,
    input [31:0] \input_data_bus_0625_wide_signal ,
    input [31:0] \input_data_bus_0626_wide_signal ,
    input [31:0] \input_data_bus_0627_wide_signal ,
    input [31:0] \input_data_bus_0628_wide_signal ,
    input [31:0] \input_data_bus_0629_wide_signal ,
    input [31:0] \input_data_bus_0630_wide_signal ,
    input [31:0] \input_data_bus_0631_wide_signal ,
    input [31:0] \input_data_bus_0632_wide_signal ,
    input [31:0] \input_data_bus_0633_wide_signal ,
    input [31:0] \input_data_bus_0634_wide_signal ,
    input [31:0] \input_data_bus_0635_wide_signal ,
    input [31:0] \input_data_bus_0636_wide_signal ,
    input [31:0] \input_data_bus_0637_wide_signal ,
    input [31:0] \input_data_bus_0638_wide_signal ,
    input [31:0] \input_data_bus_0639_wide_signal ,
    input [31:0] \input_data_bus_0640_wide_signal ,
    input [31:0] \input_data_bus_0641_wide_signal ,
    input [31:0] \input_data_bus_0642_wide_signal ,
    input [31:0] \input_data_bus_0643_wide_signal ,
    input [31:0] \input_data_bus_0644_wide_signal ,
    input [31:0] \input_data_bus_0645_wide_signal ,
    input [31:0] \input_data_bus_0646_wide_signal ,
    input [31:0] \input_data_bus_0647_wide_signal ,
    input [31:0] \input_data_bus_0648_wide_signal ,
    input [31:0] \input_data_bus_0649_wide_signal ,
    input [31:0] \input_data_bus_0650_wide_signal ,
    input [31:0] \input_data_bus_0651_wide_signal ,
    input [31:0] \input_data_bus_0652_wide_signal ,
    input [31:0] \input_data_bus_0653_wide_signal ,
    input [31:0] \input_data_bus_0654_wide_signal ,
    input [31:0] \input_data_bus_0655_wide_signal ,
    input [31:0] \input_data_bus_0656_wide_signal ,
    input [31:0] \input_data_bus_0657_wide_signal ,
    input [31:0] \input_data_bus_0658_wide_signal ,
    input [31:0] \input_data_bus_0659_wide_signal ,
    input [31:0] \input_data_bus_0660_wide_signal ,
    input [31:0] \input_data_bus_0661_wide_signal ,
    input [31:0] \input_data_bus_0662_wide_signal ,
    input [31:0] \input_data_bus_0663_wide_signal ,
    input [31:0] \input_data_bus_0664_wide_signal ,
    input [31:0] \input_data_bus_0665_wide_signal ,
    input [31:0] \input_data_bus_0666_wide_signal ,
    input [31:0] \input_data_bus_0667_wide_signal ,
    input [31:0] \input_data_bus_0668_wide_signal ,
    input [31:0] \input_data_bus_0669_wide_signal ,
    input [31:0] \input_data_bus_0670_wide_signal ,
    input [31:0] \input_data_bus_0671_wide_signal ,
    input [31:0] \input_data_bus_0672_wide_signal ,
    input [31:0] \input_data_bus_0673_wide_signal ,
    input [31:0] \input_data_bus_0674_wide_signal ,
    input [31:0] \input_data_bus_0675_wide_signal ,
    input [31:0] \input_data_bus_0676_wide_signal ,
    input [31:0] \input_data_bus_0677_wide_signal ,
    input [31:0] \input_data_bus_0678_wide_signal ,
    input [31:0] \input_data_bus_0679_wide_signal ,
    input [31:0] \input_data_bus_0680_wide_signal ,
    input [31:0] \input_data_bus_0681_wide_signal ,
    input [31:0] \input_data_bus_0682_wide_signal ,
    input [31:0] \input_data_bus_0683_wide_signal ,
    input [31:0] \input_data_bus_0684_wide_signal ,
    input [31:0] \input_data_bus_0685_wide_signal ,
    input [31:0] \input_data_bus_0686_wide_signal ,
    input [31:0] \input_data_bus_0687_wide_signal ,
    input [31:0] \input_data_bus_0688_wide_signal ,
    input [31:0] \input_data_bus_0689_wide_signal ,
    input [31:0] \input_data_bus_0690_wide_signal ,
    input [31:0] \input_data_bus_0691_wide_signal ,
    input [31:0] \input_data_bus_0692_wide_signal ,
    input [31:0] \input_data_bus_0693_wide_signal ,
    input [31:0] \input_data_bus_0694_wide_signal ,
    input [31:0] \input_data_bus_0695_wide_signal ,
    input [31:0] \input_data_bus_0696_wide_signal ,
    input [31:0] \input_data_bus_0697_wide_signal ,
    input [31:0] \input_data_bus_0698_wide_signal ,
    input [31:0] \input_data_bus_0699_wide_signal ,
    input [31:0] \input_data_bus_0700_wide_signal ,
    input [31:0] \input_data_bus_0701_wide_signal ,
    input [31:0] \input_data_bus_0702_wide_signal ,
    input [31:0] \input_data_bus_0703_wide_signal ,
    input [31:0] \input_data_bus_0704_wide_signal ,
    input [31:0] \input_data_bus_0705_wide_signal ,
    input [31:0] \input_data_bus_0706_wide_signal ,
    input [31:0] \input_data_bus_0707_wide_signal ,
    input [31:0] \input_data_bus_0708_wide_signal ,
    input [31:0] \input_data_bus_0709_wide_signal ,
    input [31:0] \input_data_bus_0710_wide_signal ,
    input [31:0] \input_data_bus_0711_wide_signal ,
    input [31:0] \input_data_bus_0712_wide_signal ,
    input [31:0] \input_data_bus_0713_wide_signal ,
    input [31:0] \input_data_bus_0714_wide_signal ,
    input [31:0] \input_data_bus_0715_wide_signal ,
    input [31:0] \input_data_bus_0716_wide_signal ,
    input [31:0] \input_data_bus_0717_wide_signal ,
    input [31:0] \input_data_bus_0718_wide_signal ,
    input [31:0] \input_data_bus_0719_wide_signal ,
    input [31:0] \input_data_bus_0720_wide_signal ,
    input [31:0] \input_data_bus_0721_wide_signal ,
    input [31:0] \input_data_bus_0722_wide_signal ,
    input [31:0] \input_data_bus_0723_wide_signal ,
    input [31:0] \input_data_bus_0724_wide_signal ,
    input [31:0] \input_data_bus_0725_wide_signal ,
    input [31:0] \input_data_bus_0726_wide_signal ,
    input [31:0] \input_data_bus_0727_wide_signal ,
    input [31:0] \input_data_bus_0728_wide_signal ,
    input [31:0] \input_data_bus_0729_wide_signal ,
    input [31:0] \input_data_bus_0730_wide_signal ,
    input [31:0] \input_data_bus_0731_wide_signal ,
    input [31:0] \input_data_bus_0732_wide_signal ,
    input [31:0] \input_data_bus_0733_wide_signal ,
    input [31:0] \input_data_bus_0734_wide_signal ,
    input [31:0] \input_data_bus_0735_wide_signal ,
    input [31:0] \input_data_bus_0736_wide_signal ,
    input [31:0] \input_data_bus_0737_wide_signal ,
    input [31:0] \input_data_bus_0738_wide_signal ,
    input [31:0] \input_data_bus_0739_wide_signal ,
    input [31:0] \input_data_bus_0740_wide_signal ,
    input [31:0] \input_data_bus_0741_wide_signal ,
    input [31:0] \input_data_bus_0742_wide_signal ,
    input [31:0] \input_data_bus_0743_wide_signal ,
    input [31:0] \input_data_bus_0744_wide_signal ,
    input [31:0] \input_data_bus_0745_wide_signal ,
    input [31:0] \input_data_bus_0746_wide_signal ,
    input [31:0] \input_data_bus_0747_wide_signal ,
    input [31:0] \input_data_bus_0748_wide_signal ,
    input [31:0] \input_data_bus_0749_wide_signal ,
    input [31:0] \input_data_bus_0750_wide_signal ,
    input [31:0] \input_data_bus_0751_wide_signal ,
    input [31:0] \input_data_bus_0752_wide_signal ,
    input [31:0] \input_data_bus_0753_wide_signal ,
    input [31:0] \input_data_bus_0754_wide_signal ,
    input [31:0] \input_data_bus_0755_wide_signal ,
    input [31:0] \input_data_bus_0756_wide_signal ,
    input [31:0] \input_data_bus_0757_wide_signal ,
    input [31:0] \input_data_bus_0758_wide_signal ,
    input [31:0] \input_data_bus_0759_wide_signal ,
    input [31:0] \input_data_bus_0760_wide_signal ,
    input [31:0] \input_data_bus_0761_wide_signal ,
    input [31:0] \input_data_bus_0762_wide_signal ,
    input [31:0] \input_data_bus_0763_wide_signal ,
    input [31:0] \input_data_bus_0764_wide_signal ,
    input [31:0] \input_data_bus_0765_wide_signal ,
    input [31:0] \input_data_bus_0766_wide_signal ,
    input [31:0] \input_data_bus_0767_wide_signal ,
    input [31:0] \input_data_bus_0768_wide_signal ,
    input [31:0] \input_data_bus_0769_wide_signal ,
    input [31:0] \input_data_bus_0770_wide_signal ,
    input [31:0] \input_data_bus_0771_wide_signal ,
    input [31:0] \input_data_bus_0772_wide_signal ,
    input [31:0] \input_data_bus_0773_wide_signal ,
    input [31:0] \input_data_bus_0774_wide_signal ,
    input [31:0] \input_data_bus_0775_wide_signal ,
    input [31:0] \input_data_bus_0776_wide_signal ,
    input [31:0] \input_data_bus_0777_wide_signal ,
    input [31:0] \input_data_bus_0778_wide_signal ,
    input [31:0] \input_data_bus_0779_wide_signal ,
    input [31:0] \input_data_bus_0780_wide_signal ,
    input [31:0] \input_data_bus_0781_wide_signal ,
    input [31:0] \input_data_bus_0782_wide_signal ,
    input [31:0] \input_data_bus_0783_wide_signal ,
    input [31:0] \input_data_bus_0784_wide_signal ,
    input [31:0] \input_data_bus_0785_wide_signal ,
    input [31:0] \input_data_bus_0786_wide_signal ,
    input [31:0] \input_data_bus_0787_wide_signal ,
    input [31:0] \input_data_bus_0788_wide_signal ,
    input [31:0] \input_data_bus_0789_wide_signal ,
    input [31:0] \input_data_bus_0790_wide_signal ,
    input [31:0] \input_data_bus_0791_wide_signal ,
    input [31:0] \input_data_bus_0792_wide_signal ,
    input [31:0] \input_data_bus_0793_wide_signal ,
    input [31:0] \input_data_bus_0794_wide_signal ,
    input [31:0] \input_data_bus_0795_wide_signal ,
    input [31:0] \input_data_bus_0796_wide_signal ,
    input [31:0] \input_data_bus_0797_wide_signal ,
    input [31:0] \input_data_bus_0798_wide_signal ,
    input [31:0] \input_data_bus_0799_wide_signal ,
    input [31:0] \input_data_bus_0800_wide_signal ,
    input [31:0] \input_data_bus_0801_wide_signal ,
    input [31:0] \input_data_bus_0802_wide_signal ,
    input [31:0] \input_data_bus_0803_wide_signal ,
    input [31:0] \input_data_bus_0804_wide_signal ,
    input [31:0] \input_data_bus_0805_wide_signal ,
    input [31:0] \input_data_bus_0806_wide_signal ,
    input [31:0] \input_data_bus_0807_wide_signal ,
    input [31:0] \input_data_bus_0808_wide_signal ,
    input [31:0] \input_data_bus_0809_wide_signal ,
    input [31:0] \input_data_bus_0810_wide_signal ,
    input [31:0] \input_data_bus_0811_wide_signal ,
    input [31:0] \input_data_bus_0812_wide_signal ,
    input [31:0] \input_data_bus_0813_wide_signal ,
    input [31:0] \input_data_bus_0814_wide_signal ,
    input [31:0] \input_data_bus_0815_wide_signal ,
    input [31:0] \input_data_bus_0816_wide_signal ,
    input [31:0] \input_data_bus_0817_wide_signal ,
    input [31:0] \input_data_bus_0818_wide_signal ,
    input [31:0] \input_data_bus_0819_wide_signal ,
    input [31:0] \input_data_bus_0820_wide_signal ,
    input [31:0] \input_data_bus_0821_wide_signal ,
    input [31:0] \input_data_bus_0822_wide_signal ,
    input [31:0] \input_data_bus_0823_wide_signal ,
    input [31:0] \input_data_bus_0824_wide_signal ,
    input [31:0] \input_data_bus_0825_wide_signal ,
    input [31:0] \input_data_bus_0826_wide_signal ,
    input [31:0] \input_data_bus_0827_wide_signal ,
    input [31:0] \input_data_bus_0828_wide_signal ,
    input [31:0] \input_data_bus_0829_wide_signal ,
    input [31:0] \input_data_bus_0830_wide_signal ,
    input [31:0] \input_data_bus_0831_wide_signal ,
    input [31:0] \input_data_bus_0832_wide_signal ,
    input [31:0] \input_data_bus_0833_wide_signal ,
    input [31:0] \input_data_bus_0834_wide_signal ,
    input [31:0] \input_data_bus_0835_wide_signal ,
    input [31:0] \input_data_bus_0836_wide_signal ,
    input [31:0] \input_data_bus_0837_wide_signal ,
    input [31:0] \input_data_bus_0838_wide_signal ,
    input [31:0] \input_data_bus_0839_wide_signal ,
    input [31:0] \input_data_bus_0840_wide_signal ,
    input [31:0] \input_data_bus_0841_wide_signal ,
    input [31:0] \input_data_bus_0842_wide_signal ,
    input [31:0] \input_data_bus_0843_wide_signal ,
    input [31:0] \input_data_bus_0844_wide_signal ,
    input [31:0] \input_data_bus_0845_wide_signal ,
    input [31:0] \input_data_bus_0846_wide_signal ,
    input [31:0] \input_data_bus_0847_wide_signal ,
    input [31:0] \input_data_bus_0848_wide_signal ,
    input [31:0] \input_data_bus_0849_wide_signal ,
    input [31:0] \input_data_bus_0850_wide_signal ,
    input [31:0] \input_data_bus_0851_wide_signal ,
    input [31:0] \input_data_bus_0852_wide_signal ,
    input [31:0] \input_data_bus_0853_wide_signal ,
    input [31:0] \input_data_bus_0854_wide_signal ,
    input [31:0] \input_data_bus_0855_wide_signal ,
    input [31:0] \input_data_bus_0856_wide_signal ,
    input [31:0] \input_data_bus_0857_wide_signal ,
    input [31:0] \input_data_bus_0858_wide_signal ,
    input [31:0] \input_data_bus_0859_wide_signal ,
    input [31:0] \input_data_bus_0860_wide_signal ,
    input [31:0] \input_data_bus_0861_wide_signal ,
    input [31:0] \input_data_bus_0862_wide_signal ,
    input [31:0] \input_data_bus_0863_wide_signal ,
    input [31:0] \input_data_bus_0864_wide_signal ,
    input [31:0] \input_data_bus_0865_wide_signal ,
    input [31:0] \input_data_bus_0866_wide_signal ,
    input [31:0] \input_data_bus_0867_wide_signal ,
    input [31:0] \input_data_bus_0868_wide_signal ,
    input [31:0] \input_data_bus_0869_wide_signal ,
    input [31:0] \input_data_bus_0870_wide_signal ,
    input [31:0] \input_data_bus_0871_wide_signal ,
    input [31:0] \input_data_bus_0872_wide_signal ,
    input [31:0] \input_data_bus_0873_wide_signal ,
    input [31:0] \input_data_bus_0874_wide_signal ,
    input [31:0] \input_data_bus_0875_wide_signal ,
    input [31:0] \input_data_bus_0876_wide_signal ,
    input [31:0] \input_data_bus_0877_wide_signal ,
    input [31:0] \input_data_bus_0878_wide_signal ,
    input [31:0] \input_data_bus_0879_wide_signal ,
    input [31:0] \input_data_bus_0880_wide_signal ,
    input [31:0] \input_data_bus_0881_wide_signal ,
    input [31:0] \input_data_bus_0882_wide_signal ,
    input [31:0] \input_data_bus_0883_wide_signal ,
    input [31:0] \input_data_bus_0884_wide_signal ,
    input [31:0] \input_data_bus_0885_wide_signal ,
    input [31:0] \input_data_bus_0886_wide_signal ,
    input [31:0] \input_data_bus_0887_wide_signal ,
    input [31:0] \input_data_bus_0888_wide_signal ,
    input [31:0] \input_data_bus_0889_wide_signal ,
    input [31:0] \input_data_bus_0890_wide_signal ,
    input [31:0] \input_data_bus_0891_wide_signal ,
    input [31:0] \input_data_bus_0892_wide_signal ,
    input [31:0] \input_data_bus_0893_wide_signal ,
    input [31:0] \input_data_bus_0894_wide_signal ,
    input [31:0] \input_data_bus_0895_wide_signal ,
    input [31:0] \input_data_bus_0896_wide_signal ,
    input [31:0] \input_data_bus_0897_wide_signal ,
    input [31:0] \input_data_bus_0898_wide_signal ,
    input [31:0] \input_data_bus_0899_wide_signal ,
    input [31:0] \input_data_bus_0900_wide_signal ,
    input [31:0] \input_data_bus_0901_wide_signal ,
    input [31:0] \input_data_bus_0902_wide_signal ,
    input [31:0] \input_data_bus_0903_wide_signal ,
    input [31:0] \input_data_bus_0904_wide_signal ,
    input [31:0] \input_data_bus_0905_wide_signal ,
    input [31:0] \input_data_bus_0906_wide_signal ,
    input [31:0] \input_data_bus_0907_wide_signal ,
    input [31:0] \input_data_bus_0908_wide_signal ,
    input [31:0] \input_data_bus_0909_wide_signal ,
    input [31:0] \input_data_bus_0910_wide_signal ,
    input [31:0] \input_data_bus_0911_wide_signal ,
    input [31:0] \input_data_bus_0912_wide_signal ,
    input [31:0] \input_data_bus_0913_wide_signal ,
    input [31:0] \input_data_bus_0914_wide_signal ,
    input [31:0] \input_data_bus_0915_wide_signal ,
    input [31:0] \input_data_bus_0916_wide_signal ,
    input [31:0] \input_data_bus_0917_wide_signal ,
    input [31:0] \input_data_bus_0918_wide_signal ,
    input [31:0] \input_data_bus_0919_wide_signal ,
    input [31:0] \input_data_bus_0920_wide_signal ,
    input [31:0] \input_data_bus_0921_wide_signal ,
    input [31:0] \input_data_bus_0922_wide_signal ,
    input [31:0] \input_data_bus_0923_wide_signal ,
    input [31:0] \input_data_bus_0924_wide_signal ,
    input [31:0] \input_data_bus_0925_wide_signal ,
    input [31:0] \input_data_bus_0926_wide_signal ,
    input [31:0] \input_data_bus_0927_wide_signal ,
    input [31:0] \input_data_bus_0928_wide_signal ,
    input [31:0] \input_data_bus_0929_wide_signal ,
    input [31:0] \input_data_bus_0930_wide_signal ,
    input [31:0] \input_data_bus_0931_wide_signal ,
    input [31:0] \input_data_bus_0932_wide_signal ,
    input [31:0] \input_data_bus_0933_wide_signal ,
    input [31:0] \input_data_bus_0934_wide_signal ,
    input [31:0] \input_data_bus_0935_wide_signal ,
    input [31:0] \input_data_bus_0936_wide_signal ,
    input [31:0] \input_data_bus_0937_wide_signal ,
    input [31:0] \input_data_bus_0938_wide_signal ,
    input [31:0] \input_data_bus_0939_wide_signal ,
    input [31:0] \input_data_bus_0940_wide_signal ,
    input [31:0] \input_data_bus_0941_wide_signal ,
    input [31:0] \input_data_bus_0942_wide_signal ,
    input [31:0] \input_data_bus_0943_wide_signal ,
    input [31:0] \input_data_bus_0944_wide_signal ,
    input [31:0] \input_data_bus_0945_wide_signal ,
    input [31:0] \input_data_bus_0946_wide_signal ,
    input [31:0] \input_data_bus_0947_wide_signal ,
    input [31:0] \input_data_bus_0948_wide_signal ,
    input [31:0] \input_data_bus_0949_wide_signal ,
    input [31:0] \input_data_bus_0950_wide_signal ,
    input [31:0] \input_data_bus_0951_wide_signal ,
    input [31:0] \input_data_bus_0952_wide_signal ,
    input [31:0] \input_data_bus_0953_wide_signal ,
    input [31:0] \input_data_bus_0954_wide_signal ,
    input [31:0] \input_data_bus_0955_wide_signal ,
    input [31:0] \input_data_bus_0956_wide_signal ,
    input [31:0] \input_data_bus_0957_wide_signal ,
    input [31:0] \input_data_bus_0958_wide_signal ,
    input [31:0] \input_data_bus_0959_wide_signal ,
    input [31:0] \input_data_bus_0960_wide_signal ,
    input [31:0] \input_data_bus_0961_wide_signal ,
    input [31:0] \input_data_bus_0962_wide_signal ,
    input [31:0] \input_data_bus_0963_wide_signal ,
    input [31:0] \input_data_bus_0964_wide_signal ,
    input [31:0] \input_data_bus_0965_wide_signal ,
    input [31:0] \input_data_bus_0966_wide_signal ,
    input [31:0] \input_data_bus_0967_wide_signal ,
    input [31:0] \input_data_bus_0968_wide_signal ,
    input [31:0] \input_data_bus_0969_wide_signal ,
    input [31:0] \input_data_bus_0970_wide_signal ,
    input [31:0] \input_data_bus_0971_wide_signal ,
    input [31:0] \input_data_bus_0972_wide_signal ,
    input [31:0] \input_data_bus_0973_wide_signal ,
    input [31:0] \input_data_bus_0974_wide_signal ,
    input [31:0] \input_data_bus_0975_wide_signal ,
    input [31:0] \input_data_bus_0976_wide_signal ,
    input [31:0] \input_data_bus_0977_wide_signal ,
    input [31:0] \input_data_bus_0978_wide_signal ,
    input [31:0] \input_data_bus_0979_wide_signal ,
    input [31:0] \input_data_bus_0980_wide_signal ,
    input [31:0] \input_data_bus_0981_wide_signal ,
    input [31:0] \input_data_bus_0982_wide_signal ,
    input [31:0] \input_data_bus_0983_wide_signal ,
    input [31:0] \input_data_bus_0984_wide_signal ,
    input [31:0] \input_data_bus_0985_wide_signal ,
    input [31:0] \input_data_bus_0986_wide_signal ,
    input [31:0] \input_data_bus_0987_wide_signal ,
    input [31:0] \input_data_bus_0988_wide_signal ,
    input [31:0] \input_data_bus_0989_wide_signal ,
    input [31:0] \input_data_bus_0990_wide_signal ,
    input [31:0] \input_data_bus_0991_wide_signal ,
    input [31:0] \input_data_bus_0992_wide_signal ,
    input [31:0] \input_data_bus_0993_wide_signal ,
    input [31:0] \input_data_bus_0994_wide_signal ,
    input [31:0] \input_data_bus_0995_wide_signal ,
    input [31:0] \input_data_bus_0996_wide_signal ,
    input [31:0] \input_data_bus_0997_wide_signal ,
    input [31:0] \input_data_bus_0998_wide_signal ,
    input [31:0] \input_data_bus_0999_wide_signal ,
    output reg [31:0] \output_data_bus_0000_wide_signal ,
    output reg [31:0] \output_data_bus_0001_wide_signal ,
    output reg [31:0] \output_data_bus_0002_wide_signal ,
    output reg [31:0] \output_data_bus_0003_wide_signal ,
    output reg [31:0] \output_data_bus_0004_wide_signal ,
    output reg [31:0] \output_data_bus_0005_wide_signal ,
    output reg [31:0] \output_data_bus_0006_wide_signal ,
    output reg [31:0] \output_data_bus_0007_wide_signal ,
    output reg [31:0] \output_data_bus_0008_wide_signal ,
    output reg [31:0] \output_data_bus_0009_wide_signal ,
    output reg [31:0] \output_data_bus_0010_wide_signal ,
    output reg [31:0] \output_data_bus_0011_wide_signal ,
    output reg [31:0] \output_data_bus_0012_wide_signal ,
    output reg [31:0] \output_data_bus_0013_wide_signal ,
    output reg [31:0] \output_data_bus_0014_wide_signal ,
    output reg [31:0] \output_data_bus_0015_wide_signal ,
    output reg [31:0] \output_data_bus_0016_wide_signal ,
    output reg [31:0] \output_data_bus_0017_wide_signal ,
    output reg [31:0] \output_data_bus_0018_wide_signal ,
    output reg [31:0] \output_data_bus_0019_wide_signal ,
    output reg [31:0] \output_data_bus_0020_wide_signal ,
    output reg [31:0] \output_data_bus_0021_wide_signal ,
    output reg [31:0] \output_data_bus_0022_wide_signal ,
    output reg [31:0] \output_data_bus_0023_wide_signal ,
    output reg [31:0] \output_data_bus_0024_wide_signal ,
    output reg [31:0] \output_data_bus_0025_wide_signal ,
    output reg [31:0] \output_data_bus_0026_wide_signal ,
    output reg [31:0] \output_data_bus_0027_wide_signal ,
    output reg [31:0] \output_data_bus_0028_wide_signal ,
    output reg [31:0] \output_data_bus_0029_wide_signal ,
    output reg [31:0] \output_data_bus_0030_wide_signal ,
    output reg [31:0] \output_data_bus_0031_wide_signal ,
    output reg [31:0] \output_data_bus_0032_wide_signal ,
    output reg [31:0] \output_data_bus_0033_wide_signal ,
    output reg [31:0] \output_data_bus_0034_wide_signal ,
    output reg [31:0] \output_data_bus_0035_wide_signal ,
    output reg [31:0] \output_data_bus_0036_wide_signal ,
    output reg [31:0] \output_data_bus_0037_wide_signal ,
    output reg [31:0] \output_data_bus_0038_wide_signal ,
    output reg [31:0] \output_data_bus_0039_wide_signal ,
    output reg [31:0] \output_data_bus_0040_wide_signal ,
    output reg [31:0] \output_data_bus_0041_wide_signal ,
    output reg [31:0] \output_data_bus_0042_wide_signal ,
    output reg [31:0] \output_data_bus_0043_wide_signal ,
    output reg [31:0] \output_data_bus_0044_wide_signal ,
    output reg [31:0] \output_data_bus_0045_wide_signal ,
    output reg [31:0] \output_data_bus_0046_wide_signal ,
    output reg [31:0] \output_data_bus_0047_wide_signal ,
    output reg [31:0] \output_data_bus_0048_wide_signal ,
    output reg [31:0] \output_data_bus_0049_wide_signal ,
    output reg [31:0] \output_data_bus_0050_wide_signal ,
    output reg [31:0] \output_data_bus_0051_wide_signal ,
    output reg [31:0] \output_data_bus_0052_wide_signal ,
    output reg [31:0] \output_data_bus_0053_wide_signal ,
    output reg [31:0] \output_data_bus_0054_wide_signal ,
    output reg [31:0] \output_data_bus_0055_wide_signal ,
    output reg [31:0] \output_data_bus_0056_wide_signal ,
    output reg [31:0] \output_data_bus_0057_wide_signal ,
    output reg [31:0] \output_data_bus_0058_wide_signal ,
    output reg [31:0] \output_data_bus_0059_wide_signal ,
    output reg [31:0] \output_data_bus_0060_wide_signal ,
    output reg [31:0] \output_data_bus_0061_wide_signal ,
    output reg [31:0] \output_data_bus_0062_wide_signal ,
    output reg [31:0] \output_data_bus_0063_wide_signal ,
    output reg [31:0] \output_data_bus_0064_wide_signal ,
    output reg [31:0] \output_data_bus_0065_wide_signal ,
    output reg [31:0] \output_data_bus_0066_wide_signal ,
    output reg [31:0] \output_data_bus_0067_wide_signal ,
    output reg [31:0] \output_data_bus_0068_wide_signal ,
    output reg [31:0] \output_data_bus_0069_wide_signal ,
    output reg [31:0] \output_data_bus_0070_wide_signal ,
    output reg [31:0] \output_data_bus_0071_wide_signal ,
    output reg [31:0] \output_data_bus_0072_wide_signal ,
    output reg [31:0] \output_data_bus_0073_wide_signal ,
    output reg [31:0] \output_data_bus_0074_wide_signal ,
    output reg [31:0] \output_data_bus_0075_wide_signal ,
    output reg [31:0] \output_data_bus_0076_wide_signal ,
    output reg [31:0] \output_data_bus_0077_wide_signal ,
    output reg [31:0] \output_data_bus_0078_wide_signal ,
    output reg [31:0] \output_data_bus_0079_wide_signal ,
    output reg [31:0] \output_data_bus_0080_wide_signal ,
    output reg [31:0] \output_data_bus_0081_wide_signal ,
    output reg [31:0] \output_data_bus_0082_wide_signal ,
    output reg [31:0] \output_data_bus_0083_wide_signal ,
    output reg [31:0] \output_data_bus_0084_wide_signal ,
    output reg [31:0] \output_data_bus_0085_wide_signal ,
    output reg [31:0] \output_data_bus_0086_wide_signal ,
    output reg [31:0] \output_data_bus_0087_wide_signal ,
    output reg [31:0] \output_data_bus_0088_wide_signal ,
    output reg [31:0] \output_data_bus_0089_wide_signal ,
    output reg [31:0] \output_data_bus_0090_wide_signal ,
    output reg [31:0] \output_data_bus_0091_wide_signal ,
    output reg [31:0] \output_data_bus_0092_wide_signal ,
    output reg [31:0] \output_data_bus_0093_wide_signal ,
    output reg [31:0] \output_data_bus_0094_wide_signal ,
    output reg [31:0] \output_data_bus_0095_wide_signal ,
    output reg [31:0] \output_data_bus_0096_wide_signal ,
    output reg [31:0] \output_data_bus_0097_wide_signal ,
    output reg [31:0] \output_data_bus_0098_wide_signal ,
    output reg [31:0] \output_data_bus_0099_wide_signal ,
    output reg [31:0] \output_data_bus_0100_wide_signal ,
    output reg [31:0] \output_data_bus_0101_wide_signal ,
    output reg [31:0] \output_data_bus_0102_wide_signal ,
    output reg [31:0] \output_data_bus_0103_wide_signal ,
    output reg [31:0] \output_data_bus_0104_wide_signal ,
    output reg [31:0] \output_data_bus_0105_wide_signal ,
    output reg [31:0] \output_data_bus_0106_wide_signal ,
    output reg [31:0] \output_data_bus_0107_wide_signal ,
    output reg [31:0] \output_data_bus_0108_wide_signal ,
    output reg [31:0] \output_data_bus_0109_wide_signal ,
    output reg [31:0] \output_data_bus_0110_wide_signal ,
    output reg [31:0] \output_data_bus_0111_wide_signal ,
    output reg [31:0] \output_data_bus_0112_wide_signal ,
    output reg [31:0] \output_data_bus_0113_wide_signal ,
    output reg [31:0] \output_data_bus_0114_wide_signal ,
    output reg [31:0] \output_data_bus_0115_wide_signal ,
    output reg [31:0] \output_data_bus_0116_wide_signal ,
    output reg [31:0] \output_data_bus_0117_wide_signal ,
    output reg [31:0] \output_data_bus_0118_wide_signal ,
    output reg [31:0] \output_data_bus_0119_wide_signal ,
    output reg [31:0] \output_data_bus_0120_wide_signal ,
    output reg [31:0] \output_data_bus_0121_wide_signal ,
    output reg [31:0] \output_data_bus_0122_wide_signal ,
    output reg [31:0] \output_data_bus_0123_wide_signal ,
    output reg [31:0] \output_data_bus_0124_wide_signal ,
    output reg [31:0] \output_data_bus_0125_wide_signal ,
    output reg [31:0] \output_data_bus_0126_wide_signal ,
    output reg [31:0] \output_data_bus_0127_wide_signal ,
    output reg [31:0] \output_data_bus_0128_wide_signal ,
    output reg [31:0] \output_data_bus_0129_wide_signal ,
    output reg [31:0] \output_data_bus_0130_wide_signal ,
    output reg [31:0] \output_data_bus_0131_wide_signal ,
    output reg [31:0] \output_data_bus_0132_wide_signal ,
    output reg [31:0] \output_data_bus_0133_wide_signal ,
    output reg [31:0] \output_data_bus_0134_wide_signal ,
    output reg [31:0] \output_data_bus_0135_wide_signal ,
    output reg [31:0] \output_data_bus_0136_wide_signal ,
    output reg [31:0] \output_data_bus_0137_wide_signal ,
    output reg [31:0] \output_data_bus_0138_wide_signal ,
    output reg [31:0] \output_data_bus_0139_wide_signal ,
    output reg [31:0] \output_data_bus_0140_wide_signal ,
    output reg [31:0] \output_data_bus_0141_wide_signal ,
    output reg [31:0] \output_data_bus_0142_wide_signal ,
    output reg [31:0] \output_data_bus_0143_wide_signal ,
    output reg [31:0] \output_data_bus_0144_wide_signal ,
    output reg [31:0] \output_data_bus_0145_wide_signal ,
    output reg [31:0] \output_data_bus_0146_wide_signal ,
    output reg [31:0] \output_data_bus_0147_wide_signal ,
    output reg [31:0] \output_data_bus_0148_wide_signal ,
    output reg [31:0] \output_data_bus_0149_wide_signal ,
    output reg [31:0] \output_data_bus_0150_wide_signal ,
    output reg [31:0] \output_data_bus_0151_wide_signal ,
    output reg [31:0] \output_data_bus_0152_wide_signal ,
    output reg [31:0] \output_data_bus_0153_wide_signal ,
    output reg [31:0] \output_data_bus_0154_wide_signal ,
    output reg [31:0] \output_data_bus_0155_wide_signal ,
    output reg [31:0] \output_data_bus_0156_wide_signal ,
    output reg [31:0] \output_data_bus_0157_wide_signal ,
    output reg [31:0] \output_data_bus_0158_wide_signal ,
    output reg [31:0] \output_data_bus_0159_wide_signal ,
    output reg [31:0] \output_data_bus_0160_wide_signal ,
    output reg [31:0] \output_data_bus_0161_wide_signal ,
    output reg [31:0] \output_data_bus_0162_wide_signal ,
    output reg [31:0] \output_data_bus_0163_wide_signal ,
    output reg [31:0] \output_data_bus_0164_wide_signal ,
    output reg [31:0] \output_data_bus_0165_wide_signal ,
    output reg [31:0] \output_data_bus_0166_wide_signal ,
    output reg [31:0] \output_data_bus_0167_wide_signal ,
    output reg [31:0] \output_data_bus_0168_wide_signal ,
    output reg [31:0] \output_data_bus_0169_wide_signal ,
    output reg [31:0] \output_data_bus_0170_wide_signal ,
    output reg [31:0] \output_data_bus_0171_wide_signal ,
    output reg [31:0] \output_data_bus_0172_wide_signal ,
    output reg [31:0] \output_data_bus_0173_wide_signal ,
    output reg [31:0] \output_data_bus_0174_wide_signal ,
    output reg [31:0] \output_data_bus_0175_wide_signal ,
    output reg [31:0] \output_data_bus_0176_wide_signal ,
    output reg [31:0] \output_data_bus_0177_wide_signal ,
    output reg [31:0] \output_data_bus_0178_wide_signal ,
    output reg [31:0] \output_data_bus_0179_wide_signal ,
    output reg [31:0] \output_data_bus_0180_wide_signal ,
    output reg [31:0] \output_data_bus_0181_wide_signal ,
    output reg [31:0] \output_data_bus_0182_wide_signal ,
    output reg [31:0] \output_data_bus_0183_wide_signal ,
    output reg [31:0] \output_data_bus_0184_wide_signal ,
    output reg [31:0] \output_data_bus_0185_wide_signal ,
    output reg [31:0] \output_data_bus_0186_wide_signal ,
    output reg [31:0] \output_data_bus_0187_wide_signal ,
    output reg [31:0] \output_data_bus_0188_wide_signal ,
    output reg [31:0] \output_data_bus_0189_wide_signal ,
    output reg [31:0] \output_data_bus_0190_wide_signal ,
    output reg [31:0] \output_data_bus_0191_wide_signal ,
    output reg [31:0] \output_data_bus_0192_wide_signal ,
    output reg [31:0] \output_data_bus_0193_wide_signal ,
    output reg [31:0] \output_data_bus_0194_wide_signal ,
    output reg [31:0] \output_data_bus_0195_wide_signal ,
    output reg [31:0] \output_data_bus_0196_wide_signal ,
    output reg [31:0] \output_data_bus_0197_wide_signal ,
    output reg [31:0] \output_data_bus_0198_wide_signal ,
    output reg [31:0] \output_data_bus_0199_wide_signal ,
    output reg [31:0] \output_data_bus_0200_wide_signal ,
    output reg [31:0] \output_data_bus_0201_wide_signal ,
    output reg [31:0] \output_data_bus_0202_wide_signal ,
    output reg [31:0] \output_data_bus_0203_wide_signal ,
    output reg [31:0] \output_data_bus_0204_wide_signal ,
    output reg [31:0] \output_data_bus_0205_wide_signal ,
    output reg [31:0] \output_data_bus_0206_wide_signal ,
    output reg [31:0] \output_data_bus_0207_wide_signal ,
    output reg [31:0] \output_data_bus_0208_wide_signal ,
    output reg [31:0] \output_data_bus_0209_wide_signal ,
    output reg [31:0] \output_data_bus_0210_wide_signal ,
    output reg [31:0] \output_data_bus_0211_wide_signal ,
    output reg [31:0] \output_data_bus_0212_wide_signal ,
    output reg [31:0] \output_data_bus_0213_wide_signal ,
    output reg [31:0] \output_data_bus_0214_wide_signal ,
    output reg [31:0] \output_data_bus_0215_wide_signal ,
    output reg [31:0] \output_data_bus_0216_wide_signal ,
    output reg [31:0] \output_data_bus_0217_wide_signal ,
    output reg [31:0] \output_data_bus_0218_wide_signal ,
    output reg [31:0] \output_data_bus_0219_wide_signal ,
    output reg [31:0] \output_data_bus_0220_wide_signal ,
    output reg [31:0] \output_data_bus_0221_wide_signal ,
    output reg [31:0] \output_data_bus_0222_wide_signal ,
    output reg [31:0] \output_data_bus_0223_wide_signal ,
    output reg [31:0] \output_data_bus_0224_wide_signal ,
    output reg [31:0] \output_data_bus_0225_wide_signal ,
    output reg [31:0] \output_data_bus_0226_wide_signal ,
    output reg [31:0] \output_data_bus_0227_wide_signal ,
    output reg [31:0] \output_data_bus_0228_wide_signal ,
    output reg [31:0] \output_data_bus_0229_wide_signal ,
    output reg [31:0] \output_data_bus_0230_wide_signal ,
    output reg [31:0] \output_data_bus_0231_wide_signal ,
    output reg [31:0] \output_data_bus_0232_wide_signal ,
    output reg [31:0] \output_data_bus_0233_wide_signal ,
    output reg [31:0] \output_data_bus_0234_wide_signal ,
    output reg [31:0] \output_data_bus_0235_wide_signal ,
    output reg [31:0] \output_data_bus_0236_wide_signal ,
    output reg [31:0] \output_data_bus_0237_wide_signal ,
    output reg [31:0] \output_data_bus_0238_wide_signal ,
    output reg [31:0] \output_data_bus_0239_wide_signal ,
    output reg [31:0] \output_data_bus_0240_wide_signal ,
    output reg [31:0] \output_data_bus_0241_wide_signal ,
    output reg [31:0] \output_data_bus_0242_wide_signal ,
    output reg [31:0] \output_data_bus_0243_wide_signal ,
    output reg [31:0] \output_data_bus_0244_wide_signal ,
    output reg [31:0] \output_data_bus_0245_wide_signal ,
    output reg [31:0] \output_data_bus_0246_wide_signal ,
    output reg [31:0] \output_data_bus_0247_wide_signal ,
    output reg [31:0] \output_data_bus_0248_wide_signal ,
    output reg [31:0] \output_data_bus_0249_wide_signal ,
    output reg [31:0] \output_data_bus_0250_wide_signal ,
    output reg [31:0] \output_data_bus_0251_wide_signal ,
    output reg [31:0] \output_data_bus_0252_wide_signal ,
    output reg [31:0] \output_data_bus_0253_wide_signal ,
    output reg [31:0] \output_data_bus_0254_wide_signal ,
    output reg [31:0] \output_data_bus_0255_wide_signal ,
    output reg [31:0] \output_data_bus_0256_wide_signal ,
    output reg [31:0] \output_data_bus_0257_wide_signal ,
    output reg [31:0] \output_data_bus_0258_wide_signal ,
    output reg [31:0] \output_data_bus_0259_wide_signal ,
    output reg [31:0] \output_data_bus_0260_wide_signal ,
    output reg [31:0] \output_data_bus_0261_wide_signal ,
    output reg [31:0] \output_data_bus_0262_wide_signal ,
    output reg [31:0] \output_data_bus_0263_wide_signal ,
    output reg [31:0] \output_data_bus_0264_wide_signal ,
    output reg [31:0] \output_data_bus_0265_wide_signal ,
    output reg [31:0] \output_data_bus_0266_wide_signal ,
    output reg [31:0] \output_data_bus_0267_wide_signal ,
    output reg [31:0] \output_data_bus_0268_wide_signal ,
    output reg [31:0] \output_data_bus_0269_wide_signal ,
    output reg [31:0] \output_data_bus_0270_wide_signal ,
    output reg [31:0] \output_data_bus_0271_wide_signal ,
    output reg [31:0] \output_data_bus_0272_wide_signal ,
    output reg [31:0] \output_data_bus_0273_wide_signal ,
    output reg [31:0] \output_data_bus_0274_wide_signal ,
    output reg [31:0] \output_data_bus_0275_wide_signal ,
    output reg [31:0] \output_data_bus_0276_wide_signal ,
    output reg [31:0] \output_data_bus_0277_wide_signal ,
    output reg [31:0] \output_data_bus_0278_wide_signal ,
    output reg [31:0] \output_data_bus_0279_wide_signal ,
    output reg [31:0] \output_data_bus_0280_wide_signal ,
    output reg [31:0] \output_data_bus_0281_wide_signal ,
    output reg [31:0] \output_data_bus_0282_wide_signal ,
    output reg [31:0] \output_data_bus_0283_wide_signal ,
    output reg [31:0] \output_data_bus_0284_wide_signal ,
    output reg [31:0] \output_data_bus_0285_wide_signal ,
    output reg [31:0] \output_data_bus_0286_wide_signal ,
    output reg [31:0] \output_data_bus_0287_wide_signal ,
    output reg [31:0] \output_data_bus_0288_wide_signal ,
    output reg [31:0] \output_data_bus_0289_wide_signal ,
    output reg [31:0] \output_data_bus_0290_wide_signal ,
    output reg [31:0] \output_data_bus_0291_wide_signal ,
    output reg [31:0] \output_data_bus_0292_wide_signal ,
    output reg [31:0] \output_data_bus_0293_wide_signal ,
    output reg [31:0] \output_data_bus_0294_wide_signal ,
    output reg [31:0] \output_data_bus_0295_wide_signal ,
    output reg [31:0] \output_data_bus_0296_wide_signal ,
    output reg [31:0] \output_data_bus_0297_wide_signal ,
    output reg [31:0] \output_data_bus_0298_wide_signal ,
    output reg [31:0] \output_data_bus_0299_wide_signal ,
    output reg [31:0] \output_data_bus_0300_wide_signal ,
    output reg [31:0] \output_data_bus_0301_wide_signal ,
    output reg [31:0] \output_data_bus_0302_wide_signal ,
    output reg [31:0] \output_data_bus_0303_wide_signal ,
    output reg [31:0] \output_data_bus_0304_wide_signal ,
    output reg [31:0] \output_data_bus_0305_wide_signal ,
    output reg [31:0] \output_data_bus_0306_wide_signal ,
    output reg [31:0] \output_data_bus_0307_wide_signal ,
    output reg [31:0] \output_data_bus_0308_wide_signal ,
    output reg [31:0] \output_data_bus_0309_wide_signal ,
    output reg [31:0] \output_data_bus_0310_wide_signal ,
    output reg [31:0] \output_data_bus_0311_wide_signal ,
    output reg [31:0] \output_data_bus_0312_wide_signal ,
    output reg [31:0] \output_data_bus_0313_wide_signal ,
    output reg [31:0] \output_data_bus_0314_wide_signal ,
    output reg [31:0] \output_data_bus_0315_wide_signal ,
    output reg [31:0] \output_data_bus_0316_wide_signal ,
    output reg [31:0] \output_data_bus_0317_wide_signal ,
    output reg [31:0] \output_data_bus_0318_wide_signal ,
    output reg [31:0] \output_data_bus_0319_wide_signal ,
    output reg [31:0] \output_data_bus_0320_wide_signal ,
    output reg [31:0] \output_data_bus_0321_wide_signal ,
    output reg [31:0] \output_data_bus_0322_wide_signal ,
    output reg [31:0] \output_data_bus_0323_wide_signal ,
    output reg [31:0] \output_data_bus_0324_wide_signal ,
    output reg [31:0] \output_data_bus_0325_wide_signal ,
    output reg [31:0] \output_data_bus_0326_wide_signal ,
    output reg [31:0] \output_data_bus_0327_wide_signal ,
    output reg [31:0] \output_data_bus_0328_wide_signal ,
    output reg [31:0] \output_data_bus_0329_wide_signal ,
    output reg [31:0] \output_data_bus_0330_wide_signal ,
    output reg [31:0] \output_data_bus_0331_wide_signal ,
    output reg [31:0] \output_data_bus_0332_wide_signal ,
    output reg [31:0] \output_data_bus_0333_wide_signal ,
    output reg [31:0] \output_data_bus_0334_wide_signal ,
    output reg [31:0] \output_data_bus_0335_wide_signal ,
    output reg [31:0] \output_data_bus_0336_wide_signal ,
    output reg [31:0] \output_data_bus_0337_wide_signal ,
    output reg [31:0] \output_data_bus_0338_wide_signal ,
    output reg [31:0] \output_data_bus_0339_wide_signal ,
    output reg [31:0] \output_data_bus_0340_wide_signal ,
    output reg [31:0] \output_data_bus_0341_wide_signal ,
    output reg [31:0] \output_data_bus_0342_wide_signal ,
    output reg [31:0] \output_data_bus_0343_wide_signal ,
    output reg [31:0] \output_data_bus_0344_wide_signal ,
    output reg [31:0] \output_data_bus_0345_wide_signal ,
    output reg [31:0] \output_data_bus_0346_wide_signal ,
    output reg [31:0] \output_data_bus_0347_wide_signal ,
    output reg [31:0] \output_data_bus_0348_wide_signal ,
    output reg [31:0] \output_data_bus_0349_wide_signal ,
    output reg [31:0] \output_data_bus_0350_wide_signal ,
    output reg [31:0] \output_data_bus_0351_wide_signal ,
    output reg [31:0] \output_data_bus_0352_wide_signal ,
    output reg [31:0] \output_data_bus_0353_wide_signal ,
    output reg [31:0] \output_data_bus_0354_wide_signal ,
    output reg [31:0] \output_data_bus_0355_wide_signal ,
    output reg [31:0] \output_data_bus_0356_wide_signal ,
    output reg [31:0] \output_data_bus_0357_wide_signal ,
    output reg [31:0] \output_data_bus_0358_wide_signal ,
    output reg [31:0] \output_data_bus_0359_wide_signal ,
    output reg [31:0] \output_data_bus_0360_wide_signal ,
    output reg [31:0] \output_data_bus_0361_wide_signal ,
    output reg [31:0] \output_data_bus_0362_wide_signal ,
    output reg [31:0] \output_data_bus_0363_wide_signal ,
    output reg [31:0] \output_data_bus_0364_wide_signal ,
    output reg [31:0] \output_data_bus_0365_wide_signal ,
    output reg [31:0] \output_data_bus_0366_wide_signal ,
    output reg [31:0] \output_data_bus_0367_wide_signal ,
    output reg [31:0] \output_data_bus_0368_wide_signal ,
    output reg [31:0] \output_data_bus_0369_wide_signal ,
    output reg [31:0] \output_data_bus_0370_wide_signal ,
    output reg [31:0] \output_data_bus_0371_wide_signal ,
    output reg [31:0] \output_data_bus_0372_wide_signal ,
    output reg [31:0] \output_data_bus_0373_wide_signal ,
    output reg [31:0] \output_data_bus_0374_wide_signal ,
    output reg [31:0] \output_data_bus_0375_wide_signal ,
    output reg [31:0] \output_data_bus_0376_wide_signal ,
    output reg [31:0] \output_data_bus_0377_wide_signal ,
    output reg [31:0] \output_data_bus_0378_wide_signal ,
    output reg [31:0] \output_data_bus_0379_wide_signal ,
    output reg [31:0] \output_data_bus_0380_wide_signal ,
    output reg [31:0] \output_data_bus_0381_wide_signal ,
    output reg [31:0] \output_data_bus_0382_wide_signal ,
    output reg [31:0] \output_data_bus_0383_wide_signal ,
    output reg [31:0] \output_data_bus_0384_wide_signal ,
    output reg [31:0] \output_data_bus_0385_wide_signal ,
    output reg [31:0] \output_data_bus_0386_wide_signal ,
    output reg [31:0] \output_data_bus_0387_wide_signal ,
    output reg [31:0] \output_data_bus_0388_wide_signal ,
    output reg [31:0] \output_data_bus_0389_wide_signal ,
    output reg [31:0] \output_data_bus_0390_wide_signal ,
    output reg [31:0] \output_data_bus_0391_wide_signal ,
    output reg [31:0] \output_data_bus_0392_wide_signal ,
    output reg [31:0] \output_data_bus_0393_wide_signal ,
    output reg [31:0] \output_data_bus_0394_wide_signal ,
    output reg [31:0] \output_data_bus_0395_wide_signal ,
    output reg [31:0] \output_data_bus_0396_wide_signal ,
    output reg [31:0] \output_data_bus_0397_wide_signal ,
    output reg [31:0] \output_data_bus_0398_wide_signal ,
    output reg [31:0] \output_data_bus_0399_wide_signal ,
    output reg [31:0] \output_data_bus_0400_wide_signal ,
    output reg [31:0] \output_data_bus_0401_wide_signal ,
    output reg [31:0] \output_data_bus_0402_wide_signal ,
    output reg [31:0] \output_data_bus_0403_wide_signal ,
    output reg [31:0] \output_data_bus_0404_wide_signal ,
    output reg [31:0] \output_data_bus_0405_wide_signal ,
    output reg [31:0] \output_data_bus_0406_wide_signal ,
    output reg [31:0] \output_data_bus_0407_wide_signal ,
    output reg [31:0] \output_data_bus_0408_wide_signal ,
    output reg [31:0] \output_data_bus_0409_wide_signal ,
    output reg [31:0] \output_data_bus_0410_wide_signal ,
    output reg [31:0] \output_data_bus_0411_wide_signal ,
    output reg [31:0] \output_data_bus_0412_wide_signal ,
    output reg [31:0] \output_data_bus_0413_wide_signal ,
    output reg [31:0] \output_data_bus_0414_wide_signal ,
    output reg [31:0] \output_data_bus_0415_wide_signal ,
    output reg [31:0] \output_data_bus_0416_wide_signal ,
    output reg [31:0] \output_data_bus_0417_wide_signal ,
    output reg [31:0] \output_data_bus_0418_wide_signal ,
    output reg [31:0] \output_data_bus_0419_wide_signal ,
    output reg [31:0] \output_data_bus_0420_wide_signal ,
    output reg [31:0] \output_data_bus_0421_wide_signal ,
    output reg [31:0] \output_data_bus_0422_wide_signal ,
    output reg [31:0] \output_data_bus_0423_wide_signal ,
    output reg [31:0] \output_data_bus_0424_wide_signal ,
    output reg [31:0] \output_data_bus_0425_wide_signal ,
    output reg [31:0] \output_data_bus_0426_wide_signal ,
    output reg [31:0] \output_data_bus_0427_wide_signal ,
    output reg [31:0] \output_data_bus_0428_wide_signal ,
    output reg [31:0] \output_data_bus_0429_wide_signal ,
    output reg [31:0] \output_data_bus_0430_wide_signal ,
    output reg [31:0] \output_data_bus_0431_wide_signal ,
    output reg [31:0] \output_data_bus_0432_wide_signal ,
    output reg [31:0] \output_data_bus_0433_wide_signal ,
    output reg [31:0] \output_data_bus_0434_wide_signal ,
    output reg [31:0] \output_data_bus_0435_wide_signal ,
    output reg [31:0] \output_data_bus_0436_wide_signal ,
    output reg [31:0] \output_data_bus_0437_wide_signal ,
    output reg [31:0] \output_data_bus_0438_wide_signal ,
    output reg [31:0] \output_data_bus_0439_wide_signal ,
    output reg [31:0] \output_data_bus_0440_wide_signal ,
    output reg [31:0] \output_data_bus_0441_wide_signal ,
    output reg [31:0] \output_data_bus_0442_wide_signal ,
    output reg [31:0] \output_data_bus_0443_wide_signal ,
    output reg [31:0] \output_data_bus_0444_wide_signal ,
    output reg [31:0] \output_data_bus_0445_wide_signal ,
    output reg [31:0] \output_data_bus_0446_wide_signal ,
    output reg [31:0] \output_data_bus_0447_wide_signal ,
    output reg [31:0] \output_data_bus_0448_wide_signal ,
    output reg [31:0] \output_data_bus_0449_wide_signal ,
    output reg [31:0] \output_data_bus_0450_wide_signal ,
    output reg [31:0] \output_data_bus_0451_wide_signal ,
    output reg [31:0] \output_data_bus_0452_wide_signal ,
    output reg [31:0] \output_data_bus_0453_wide_signal ,
    output reg [31:0] \output_data_bus_0454_wide_signal ,
    output reg [31:0] \output_data_bus_0455_wide_signal ,
    output reg [31:0] \output_data_bus_0456_wide_signal ,
    output reg [31:0] \output_data_bus_0457_wide_signal ,
    output reg [31:0] \output_data_bus_0458_wide_signal ,
    output reg [31:0] \output_data_bus_0459_wide_signal ,
    output reg [31:0] \output_data_bus_0460_wide_signal ,
    output reg [31:0] \output_data_bus_0461_wide_signal ,
    output reg [31:0] \output_data_bus_0462_wide_signal ,
    output reg [31:0] \output_data_bus_0463_wide_signal ,
    output reg [31:0] \output_data_bus_0464_wide_signal ,
    output reg [31:0] \output_data_bus_0465_wide_signal ,
    output reg [31:0] \output_data_bus_0466_wide_signal ,
    output reg [31:0] \output_data_bus_0467_wide_signal ,
    output reg [31:0] \output_data_bus_0468_wide_signal ,
    output reg [31:0] \output_data_bus_0469_wide_signal ,
    output reg [31:0] \output_data_bus_0470_wide_signal ,
    output reg [31:0] \output_data_bus_0471_wide_signal ,
    output reg [31:0] \output_data_bus_0472_wide_signal ,
    output reg [31:0] \output_data_bus_0473_wide_signal ,
    output reg [31:0] \output_data_bus_0474_wide_signal ,
    output reg [31:0] \output_data_bus_0475_wide_signal ,
    output reg [31:0] \output_data_bus_0476_wide_signal ,
    output reg [31:0] \output_data_bus_0477_wide_signal ,
    output reg [31:0] \output_data_bus_0478_wide_signal ,
    output reg [31:0] \output_data_bus_0479_wide_signal ,
    output reg [31:0] \output_data_bus_0480_wide_signal ,
    output reg [31:0] \output_data_bus_0481_wide_signal ,
    output reg [31:0] \output_data_bus_0482_wide_signal ,
    output reg [31:0] \output_data_bus_0483_wide_signal ,
    output reg [31:0] \output_data_bus_0484_wide_signal ,
    output reg [31:0] \output_data_bus_0485_wide_signal ,
    output reg [31:0] \output_data_bus_0486_wide_signal ,
    output reg [31:0] \output_data_bus_0487_wide_signal ,
    output reg [31:0] \output_data_bus_0488_wide_signal ,
    output reg [31:0] \output_data_bus_0489_wide_signal ,
    output reg [31:0] \output_data_bus_0490_wide_signal ,
    output reg [31:0] \output_data_bus_0491_wide_signal ,
    output reg [31:0] \output_data_bus_0492_wide_signal ,
    output reg [31:0] \output_data_bus_0493_wide_signal ,
    output reg [31:0] \output_data_bus_0494_wide_signal ,
    output reg [31:0] \output_data_bus_0495_wide_signal ,
    output reg [31:0] \output_data_bus_0496_wide_signal ,
    output reg [31:0] \output_data_bus_0497_wide_signal ,
    output reg [31:0] \output_data_bus_0498_wide_signal ,
    output reg [31:0] \output_data_bus_0499_wide_signal ,
    output reg [31:0] \output_data_bus_0500_wide_signal ,
    output reg [31:0] \output_data_bus_0501_wide_signal ,
    output reg [31:0] \output_data_bus_0502_wide_signal ,
    output reg [31:0] \output_data_bus_0503_wide_signal ,
    output reg [31:0] \output_data_bus_0504_wide_signal ,
    output reg [31:0] \output_data_bus_0505_wide_signal ,
    output reg [31:0] \output_data_bus_0506_wide_signal ,
    output reg [31:0] \output_data_bus_0507_wide_signal ,
    output reg [31:0] \output_data_bus_0508_wide_signal ,
    output reg [31:0] \output_data_bus_0509_wide_signal ,
    output reg [31:0] \output_data_bus_0510_wide_signal ,
    output reg [31:0] \output_data_bus_0511_wide_signal ,
    output reg [31:0] \output_data_bus_0512_wide_signal ,
    output reg [31:0] \output_data_bus_0513_wide_signal ,
    output reg [31:0] \output_data_bus_0514_wide_signal ,
    output reg [31:0] \output_data_bus_0515_wide_signal ,
    output reg [31:0] \output_data_bus_0516_wide_signal ,
    output reg [31:0] \output_data_bus_0517_wide_signal ,
    output reg [31:0] \output_data_bus_0518_wide_signal ,
    output reg [31:0] \output_data_bus_0519_wide_signal ,
    output reg [31:0] \output_data_bus_0520_wide_signal ,
    output reg [31:0] \output_data_bus_0521_wide_signal ,
    output reg [31:0] \output_data_bus_0522_wide_signal ,
    output reg [31:0] \output_data_bus_0523_wide_signal ,
    output reg [31:0] \output_data_bus_0524_wide_signal ,
    output reg [31:0] \output_data_bus_0525_wide_signal ,
    output reg [31:0] \output_data_bus_0526_wide_signal ,
    output reg [31:0] \output_data_bus_0527_wide_signal ,
    output reg [31:0] \output_data_bus_0528_wide_signal ,
    output reg [31:0] \output_data_bus_0529_wide_signal ,
    output reg [31:0] \output_data_bus_0530_wide_signal ,
    output reg [31:0] \output_data_bus_0531_wide_signal ,
    output reg [31:0] \output_data_bus_0532_wide_signal ,
    output reg [31:0] \output_data_bus_0533_wide_signal ,
    output reg [31:0] \output_data_bus_0534_wide_signal ,
    output reg [31:0] \output_data_bus_0535_wide_signal ,
    output reg [31:0] \output_data_bus_0536_wide_signal ,
    output reg [31:0] \output_data_bus_0537_wide_signal ,
    output reg [31:0] \output_data_bus_0538_wide_signal ,
    output reg [31:0] \output_data_bus_0539_wide_signal ,
    output reg [31:0] \output_data_bus_0540_wide_signal ,
    output reg [31:0] \output_data_bus_0541_wide_signal ,
    output reg [31:0] \output_data_bus_0542_wide_signal ,
    output reg [31:0] \output_data_bus_0543_wide_signal ,
    output reg [31:0] \output_data_bus_0544_wide_signal ,
    output reg [31:0] \output_data_bus_0545_wide_signal ,
    output reg [31:0] \output_data_bus_0546_wide_signal ,
    output reg [31:0] \output_data_bus_0547_wide_signal ,
    output reg [31:0] \output_data_bus_0548_wide_signal ,
    output reg [31:0] \output_data_bus_0549_wide_signal ,
    output reg [31:0] \output_data_bus_0550_wide_signal ,
    output reg [31:0] \output_data_bus_0551_wide_signal ,
    output reg [31:0] \output_data_bus_0552_wide_signal ,
    output reg [31:0] \output_data_bus_0553_wide_signal ,
    output reg [31:0] \output_data_bus_0554_wide_signal ,
    output reg [31:0] \output_data_bus_0555_wide_signal ,
    output reg [31:0] \output_data_bus_0556_wide_signal ,
    output reg [31:0] \output_data_bus_0557_wide_signal ,
    output reg [31:0] \output_data_bus_0558_wide_signal ,
    output reg [31:0] \output_data_bus_0559_wide_signal ,
    output reg [31:0] \output_data_bus_0560_wide_signal ,
    output reg [31:0] \output_data_bus_0561_wide_signal ,
    output reg [31:0] \output_data_bus_0562_wide_signal ,
    output reg [31:0] \output_data_bus_0563_wide_signal ,
    output reg [31:0] \output_data_bus_0564_wide_signal ,
    output reg [31:0] \output_data_bus_0565_wide_signal ,
    output reg [31:0] \output_data_bus_0566_wide_signal ,
    output reg [31:0] \output_data_bus_0567_wide_signal ,
    output reg [31:0] \output_data_bus_0568_wide_signal ,
    output reg [31:0] \output_data_bus_0569_wide_signal ,
    output reg [31:0] \output_data_bus_0570_wide_signal ,
    output reg [31:0] \output_data_bus_0571_wide_signal ,
    output reg [31:0] \output_data_bus_0572_wide_signal ,
    output reg [31:0] \output_data_bus_0573_wide_signal ,
    output reg [31:0] \output_data_bus_0574_wide_signal ,
    output reg [31:0] \output_data_bus_0575_wide_signal ,
    output reg [31:0] \output_data_bus_0576_wide_signal ,
    output reg [31:0] \output_data_bus_0577_wide_signal ,
    output reg [31:0] \output_data_bus_0578_wide_signal ,
    output reg [31:0] \output_data_bus_0579_wide_signal ,
    output reg [31:0] \output_data_bus_0580_wide_signal ,
    output reg [31:0] \output_data_bus_0581_wide_signal ,
    output reg [31:0] \output_data_bus_0582_wide_signal ,
    output reg [31:0] \output_data_bus_0583_wide_signal ,
    output reg [31:0] \output_data_bus_0584_wide_signal ,
    output reg [31:0] \output_data_bus_0585_wide_signal ,
    output reg [31:0] \output_data_bus_0586_wide_signal ,
    output reg [31:0] \output_data_bus_0587_wide_signal ,
    output reg [31:0] \output_data_bus_0588_wide_signal ,
    output reg [31:0] \output_data_bus_0589_wide_signal ,
    output reg [31:0] \output_data_bus_0590_wide_signal ,
    output reg [31:0] \output_data_bus_0591_wide_signal ,
    output reg [31:0] \output_data_bus_0592_wide_signal ,
    output reg [31:0] \output_data_bus_0593_wide_signal ,
    output reg [31:0] \output_data_bus_0594_wide_signal ,
    output reg [31:0] \output_data_bus_0595_wide_signal ,
    output reg [31:0] \output_data_bus_0596_wide_signal ,
    output reg [31:0] \output_data_bus_0597_wide_signal ,
    output reg [31:0] \output_data_bus_0598_wide_signal ,
    output reg [31:0] \output_data_bus_0599_wide_signal ,
    output reg [31:0] \output_data_bus_0600_wide_signal ,
    output reg [31:0] \output_data_bus_0601_wide_signal ,
    output reg [31:0] \output_data_bus_0602_wide_signal ,
    output reg [31:0] \output_data_bus_0603_wide_signal ,
    output reg [31:0] \output_data_bus_0604_wide_signal ,
    output reg [31:0] \output_data_bus_0605_wide_signal ,
    output reg [31:0] \output_data_bus_0606_wide_signal ,
    output reg [31:0] \output_data_bus_0607_wide_signal ,
    output reg [31:0] \output_data_bus_0608_wide_signal ,
    output reg [31:0] \output_data_bus_0609_wide_signal ,
    output reg [31:0] \output_data_bus_0610_wide_signal ,
    output reg [31:0] \output_data_bus_0611_wide_signal ,
    output reg [31:0] \output_data_bus_0612_wide_signal ,
    output reg [31:0] \output_data_bus_0613_wide_signal ,
    output reg [31:0] \output_data_bus_0614_wide_signal ,
    output reg [31:0] \output_data_bus_0615_wide_signal ,
    output reg [31:0] \output_data_bus_0616_wide_signal ,
    output reg [31:0] \output_data_bus_0617_wide_signal ,
    output reg [31:0] \output_data_bus_0618_wide_signal ,
    output reg [31:0] \output_data_bus_0619_wide_signal ,
    output reg [31:0] \output_data_bus_0620_wide_signal ,
    output reg [31:0] \output_data_bus_0621_wide_signal ,
    output reg [31:0] \output_data_bus_0622_wide_signal ,
    output reg [31:0] \output_data_bus_0623_wide_signal ,
    output reg [31:0] \output_data_bus_0624_wide_signal ,
    output reg [31:0] \output_data_bus_0625_wide_signal ,
    output reg [31:0] \output_data_bus_0626_wide_signal ,
    output reg [31:0] \output_data_bus_0627_wide_signal ,
    output reg [31:0] \output_data_bus_0628_wide_signal ,
    output reg [31:0] \output_data_bus_0629_wide_signal ,
    output reg [31:0] \output_data_bus_0630_wide_signal ,
    output reg [31:0] \output_data_bus_0631_wide_signal ,
    output reg [31:0] \output_data_bus_0632_wide_signal ,
    output reg [31:0] \output_data_bus_0633_wide_signal ,
    output reg [31:0] \output_data_bus_0634_wide_signal ,
    output reg [31:0] \output_data_bus_0635_wide_signal ,
    output reg [31:0] \output_data_bus_0636_wide_signal ,
    output reg [31:0] \output_data_bus_0637_wide_signal ,
    output reg [31:0] \output_data_bus_0638_wide_signal ,
    output reg [31:0] \output_data_bus_0639_wide_signal ,
    output reg [31:0] \output_data_bus_0640_wide_signal ,
    output reg [31:0] \output_data_bus_0641_wide_signal ,
    output reg [31:0] \output_data_bus_0642_wide_signal ,
    output reg [31:0] \output_data_bus_0643_wide_signal ,
    output reg [31:0] \output_data_bus_0644_wide_signal ,
    output reg [31:0] \output_data_bus_0645_wide_signal ,
    output reg [31:0] \output_data_bus_0646_wide_signal ,
    output reg [31:0] \output_data_bus_0647_wide_signal ,
    output reg [31:0] \output_data_bus_0648_wide_signal ,
    output reg [31:0] \output_data_bus_0649_wide_signal ,
    output reg [31:0] \output_data_bus_0650_wide_signal ,
    output reg [31:0] \output_data_bus_0651_wide_signal ,
    output reg [31:0] \output_data_bus_0652_wide_signal ,
    output reg [31:0] \output_data_bus_0653_wide_signal ,
    output reg [31:0] \output_data_bus_0654_wide_signal ,
    output reg [31:0] \output_data_bus_0655_wide_signal ,
    output reg [31:0] \output_data_bus_0656_wide_signal ,
    output reg [31:0] \output_data_bus_0657_wide_signal ,
    output reg [31:0] \output_data_bus_0658_wide_signal ,
    output reg [31:0] \output_data_bus_0659_wide_signal ,
    output reg [31:0] \output_data_bus_0660_wide_signal ,
    output reg [31:0] \output_data_bus_0661_wide_signal ,
    output reg [31:0] \output_data_bus_0662_wide_signal ,
    output reg [31:0] \output_data_bus_0663_wide_signal ,
    output reg [31:0] \output_data_bus_0664_wide_signal ,
    output reg [31:0] \output_data_bus_0665_wide_signal ,
    output reg [31:0] \output_data_bus_0666_wide_signal ,
    output reg [31:0] \output_data_bus_0667_wide_signal ,
    output reg [31:0] \output_data_bus_0668_wide_signal ,
    output reg [31:0] \output_data_bus_0669_wide_signal ,
    output reg [31:0] \output_data_bus_0670_wide_signal ,
    output reg [31:0] \output_data_bus_0671_wide_signal ,
    output reg [31:0] \output_data_bus_0672_wide_signal ,
    output reg [31:0] \output_data_bus_0673_wide_signal ,
    output reg [31:0] \output_data_bus_0674_wide_signal ,
    output reg [31:0] \output_data_bus_0675_wide_signal ,
    output reg [31:0] \output_data_bus_0676_wide_signal ,
    output reg [31:0] \output_data_bus_0677_wide_signal ,
    output reg [31:0] \output_data_bus_0678_wide_signal ,
    output reg [31:0] \output_data_bus_0679_wide_signal ,
    output reg [31:0] \output_data_bus_0680_wide_signal ,
    output reg [31:0] \output_data_bus_0681_wide_signal ,
    output reg [31:0] \output_data_bus_0682_wide_signal ,
    output reg [31:0] \output_data_bus_0683_wide_signal ,
    output reg [31:0] \output_data_bus_0684_wide_signal ,
    output reg [31:0] \output_data_bus_0685_wide_signal ,
    output reg [31:0] \output_data_bus_0686_wide_signal ,
    output reg [31:0] \output_data_bus_0687_wide_signal ,
    output reg [31:0] \output_data_bus_0688_wide_signal ,
    output reg [31:0] \output_data_bus_0689_wide_signal ,
    output reg [31:0] \output_data_bus_0690_wide_signal ,
    output reg [31:0] \output_data_bus_0691_wide_signal ,
    output reg [31:0] \output_data_bus_0692_wide_signal ,
    output reg [31:0] \output_data_bus_0693_wide_signal ,
    output reg [31:0] \output_data_bus_0694_wide_signal ,
    output reg [31:0] \output_data_bus_0695_wide_signal ,
    output reg [31:0] \output_data_bus_0696_wide_signal ,
    output reg [31:0] \output_data_bus_0697_wide_signal ,
    output reg [31:0] \output_data_bus_0698_wide_signal ,
    output reg [31:0] \output_data_bus_0699_wide_signal ,
    output reg [31:0] \output_data_bus_0700_wide_signal ,
    output reg [31:0] \output_data_bus_0701_wide_signal ,
    output reg [31:0] \output_data_bus_0702_wide_signal ,
    output reg [31:0] \output_data_bus_0703_wide_signal ,
    output reg [31:0] \output_data_bus_0704_wide_signal ,
    output reg [31:0] \output_data_bus_0705_wide_signal ,
    output reg [31:0] \output_data_bus_0706_wide_signal ,
    output reg [31:0] \output_data_bus_0707_wide_signal ,
    output reg [31:0] \output_data_bus_0708_wide_signal ,
    output reg [31:0] \output_data_bus_0709_wide_signal ,
    output reg [31:0] \output_data_bus_0710_wide_signal ,
    output reg [31:0] \output_data_bus_0711_wide_signal ,
    output reg [31:0] \output_data_bus_0712_wide_signal ,
    output reg [31:0] \output_data_bus_0713_wide_signal ,
    output reg [31:0] \output_data_bus_0714_wide_signal ,
    output reg [31:0] \output_data_bus_0715_wide_signal ,
    output reg [31:0] \output_data_bus_0716_wide_signal ,
    output reg [31:0] \output_data_bus_0717_wide_signal ,
    output reg [31:0] \output_data_bus_0718_wide_signal ,
    output reg [31:0] \output_data_bus_0719_wide_signal ,
    output reg [31:0] \output_data_bus_0720_wide_signal ,
    output reg [31:0] \output_data_bus_0721_wide_signal ,
    output reg [31:0] \output_data_bus_0722_wide_signal ,
    output reg [31:0] \output_data_bus_0723_wide_signal ,
    output reg [31:0] \output_data_bus_0724_wide_signal ,
    output reg [31:0] \output_data_bus_0725_wide_signal ,
    output reg [31:0] \output_data_bus_0726_wide_signal ,
    output reg [31:0] \output_data_bus_0727_wide_signal ,
    output reg [31:0] \output_data_bus_0728_wide_signal ,
    output reg [31:0] \output_data_bus_0729_wide_signal ,
    output reg [31:0] \output_data_bus_0730_wide_signal ,
    output reg [31:0] \output_data_bus_0731_wide_signal ,
    output reg [31:0] \output_data_bus_0732_wide_signal ,
    output reg [31:0] \output_data_bus_0733_wide_signal ,
    output reg [31:0] \output_data_bus_0734_wide_signal ,
    output reg [31:0] \output_data_bus_0735_wide_signal ,
    output reg [31:0] \output_data_bus_0736_wide_signal ,
    output reg [31:0] \output_data_bus_0737_wide_signal ,
    output reg [31:0] \output_data_bus_0738_wide_signal ,
    output reg [31:0] \output_data_bus_0739_wide_signal ,
    output reg [31:0] \output_data_bus_0740_wide_signal ,
    output reg [31:0] \output_data_bus_0741_wide_signal ,
    output reg [31:0] \output_data_bus_0742_wide_signal ,
    output reg [31:0] \output_data_bus_0743_wide_signal ,
    output reg [31:0] \output_data_bus_0744_wide_signal ,
    output reg [31:0] \output_data_bus_0745_wide_signal ,
    output reg [31:0] \output_data_bus_0746_wide_signal ,
    output reg [31:0] \output_data_bus_0747_wide_signal ,
    output reg [31:0] \output_data_bus_0748_wide_signal ,
    output reg [31:0] \output_data_bus_0749_wide_signal ,
    output reg [31:0] \output_data_bus_0750_wide_signal ,
    output reg [31:0] \output_data_bus_0751_wide_signal ,
    output reg [31:0] \output_data_bus_0752_wide_signal ,
    output reg [31:0] \output_data_bus_0753_wide_signal ,
    output reg [31:0] \output_data_bus_0754_wide_signal ,
    output reg [31:0] \output_data_bus_0755_wide_signal ,
    output reg [31:0] \output_data_bus_0756_wide_signal ,
    output reg [31:0] \output_data_bus_0757_wide_signal ,
    output reg [31:0] \output_data_bus_0758_wide_signal ,
    output reg [31:0] \output_data_bus_0759_wide_signal ,
    output reg [31:0] \output_data_bus_0760_wide_signal ,
    output reg [31:0] \output_data_bus_0761_wide_signal ,
    output reg [31:0] \output_data_bus_0762_wide_signal ,
    output reg [31:0] \output_data_bus_0763_wide_signal ,
    output reg [31:0] \output_data_bus_0764_wide_signal ,
    output reg [31:0] \output_data_bus_0765_wide_signal ,
    output reg [31:0] \output_data_bus_0766_wide_signal ,
    output reg [31:0] \output_data_bus_0767_wide_signal ,
    output reg [31:0] \output_data_bus_0768_wide_signal ,
    output reg [31:0] \output_data_bus_0769_wide_signal ,
    output reg [31:0] \output_data_bus_0770_wide_signal ,
    output reg [31:0] \output_data_bus_0771_wide_signal ,
    output reg [31:0] \output_data_bus_0772_wide_signal ,
    output reg [31:0] \output_data_bus_0773_wide_signal ,
    output reg [31:0] \output_data_bus_0774_wide_signal ,
    output reg [31:0] \output_data_bus_0775_wide_signal ,
    output reg [31:0] \output_data_bus_0776_wide_signal ,
    output reg [31:0] \output_data_bus_0777_wide_signal ,
    output reg [31:0] \output_data_bus_0778_wide_signal ,
    output reg [31:0] \output_data_bus_0779_wide_signal ,
    output reg [31:0] \output_data_bus_0780_wide_signal ,
    output reg [31:0] \output_data_bus_0781_wide_signal ,
    output reg [31:0] \output_data_bus_0782_wide_signal ,
    output reg [31:0] \output_data_bus_0783_wide_signal ,
    output reg [31:0] \output_data_bus_0784_wide_signal ,
    output reg [31:0] \output_data_bus_0785_wide_signal ,
    output reg [31:0] \output_data_bus_0786_wide_signal ,
    output reg [31:0] \output_data_bus_0787_wide_signal ,
    output reg [31:0] \output_data_bus_0788_wide_signal ,
    output reg [31:0] \output_data_bus_0789_wide_signal ,
    output reg [31:0] \output_data_bus_0790_wide_signal ,
    output reg [31:0] \output_data_bus_0791_wide_signal ,
    output reg [31:0] \output_data_bus_0792_wide_signal ,
    output reg [31:0] \output_data_bus_0793_wide_signal ,
    output reg [31:0] \output_data_bus_0794_wide_signal ,
    output reg [31:0] \output_data_bus_0795_wide_signal ,
    output reg [31:0] \output_data_bus_0796_wide_signal ,
    output reg [31:0] \output_data_bus_0797_wide_signal ,
    output reg [31:0] \output_data_bus_0798_wide_signal ,
    output reg [31:0] \output_data_bus_0799_wide_signal ,
    output reg [31:0] \output_data_bus_0800_wide_signal ,
    output reg [31:0] \output_data_bus_0801_wide_signal ,
    output reg [31:0] \output_data_bus_0802_wide_signal ,
    output reg [31:0] \output_data_bus_0803_wide_signal ,
    output reg [31:0] \output_data_bus_0804_wide_signal ,
    output reg [31:0] \output_data_bus_0805_wide_signal ,
    output reg [31:0] \output_data_bus_0806_wide_signal ,
    output reg [31:0] \output_data_bus_0807_wide_signal ,
    output reg [31:0] \output_data_bus_0808_wide_signal ,
    output reg [31:0] \output_data_bus_0809_wide_signal ,
    output reg [31:0] \output_data_bus_0810_wide_signal ,
    output reg [31:0] \output_data_bus_0811_wide_signal ,
    output reg [31:0] \output_data_bus_0812_wide_signal ,
    output reg [31:0] \output_data_bus_0813_wide_signal ,
    output reg [31:0] \output_data_bus_0814_wide_signal ,
    output reg [31:0] \output_data_bus_0815_wide_signal ,
    output reg [31:0] \output_data_bus_0816_wide_signal ,
    output reg [31:0] \output_data_bus_0817_wide_signal ,
    output reg [31:0] \output_data_bus_0818_wide_signal ,
    output reg [31:0] \output_data_bus_0819_wide_signal ,
    output reg [31:0] \output_data_bus_0820_wide_signal ,
    output reg [31:0] \output_data_bus_0821_wide_signal ,
    output reg [31:0] \output_data_bus_0822_wide_signal ,
    output reg [31:0] \output_data_bus_0823_wide_signal ,
    output reg [31:0] \output_data_bus_0824_wide_signal ,
    output reg [31:0] \output_data_bus_0825_wide_signal ,
    output reg [31:0] \output_data_bus_0826_wide_signal ,
    output reg [31:0] \output_data_bus_0827_wide_signal ,
    output reg [31:0] \output_data_bus_0828_wide_signal ,
    output reg [31:0] \output_data_bus_0829_wide_signal ,
    output reg [31:0] \output_data_bus_0830_wide_signal ,
    output reg [31:0] \output_data_bus_0831_wide_signal ,
    output reg [31:0] \output_data_bus_0832_wide_signal ,
    output reg [31:0] \output_data_bus_0833_wide_signal ,
    output reg [31:0] \output_data_bus_0834_wide_signal ,
    output reg [31:0] \output_data_bus_0835_wide_signal ,
    output reg [31:0] \output_data_bus_0836_wide_signal ,
    output reg [31:0] \output_data_bus_0837_wide_signal ,
    output reg [31:0] \output_data_bus_0838_wide_signal ,
    output reg [31:0] \output_data_bus_0839_wide_signal ,
    output reg [31:0] \output_data_bus_0840_wide_signal ,
    output reg [31:0] \output_data_bus_0841_wide_signal ,
    output reg [31:0] \output_data_bus_0842_wide_signal ,
    output reg [31:0] \output_data_bus_0843_wide_signal ,
    output reg [31:0] \output_data_bus_0844_wide_signal ,
    output reg [31:0] \output_data_bus_0845_wide_signal ,
    output reg [31:0] \output_data_bus_0846_wide_signal ,
    output reg [31:0] \output_data_bus_0847_wide_signal ,
    output reg [31:0] \output_data_bus_0848_wide_signal ,
    output reg [31:0] \output_data_bus_0849_wide_signal ,
    output reg [31:0] \output_data_bus_0850_wide_signal ,
    output reg [31:0] \output_data_bus_0851_wide_signal ,
    output reg [31:0] \output_data_bus_0852_wide_signal ,
    output reg [31:0] \output_data_bus_0853_wide_signal ,
    output reg [31:0] \output_data_bus_0854_wide_signal ,
    output reg [31:0] \output_data_bus_0855_wide_signal ,
    output reg [31:0] \output_data_bus_0856_wide_signal ,
    output reg [31:0] \output_data_bus_0857_wide_signal ,
    output reg [31:0] \output_data_bus_0858_wide_signal ,
    output reg [31:0] \output_data_bus_0859_wide_signal ,
    output reg [31:0] \output_data_bus_0860_wide_signal ,
    output reg [31:0] \output_data_bus_0861_wide_signal ,
    output reg [31:0] \output_data_bus_0862_wide_signal ,
    output reg [31:0] \output_data_bus_0863_wide_signal ,
    output reg [31:0] \output_data_bus_0864_wide_signal ,
    output reg [31:0] \output_data_bus_0865_wide_signal ,
    output reg [31:0] \output_data_bus_0866_wide_signal ,
    output reg [31:0] \output_data_bus_0867_wide_signal ,
    output reg [31:0] \output_data_bus_0868_wide_signal ,
    output reg [31:0] \output_data_bus_0869_wide_signal ,
    output reg [31:0] \output_data_bus_0870_wide_signal ,
    output reg [31:0] \output_data_bus_0871_wide_signal ,
    output reg [31:0] \output_data_bus_0872_wide_signal ,
    output reg [31:0] \output_data_bus_0873_wide_signal ,
    output reg [31:0] \output_data_bus_0874_wide_signal ,
    output reg [31:0] \output_data_bus_0875_wide_signal ,
    output reg [31:0] \output_data_bus_0876_wide_signal ,
    output reg [31:0] \output_data_bus_0877_wide_signal ,
    output reg [31:0] \output_data_bus_0878_wide_signal ,
    output reg [31:0] \output_data_bus_0879_wide_signal ,
    output reg [31:0] \output_data_bus_0880_wide_signal ,
    output reg [31:0] \output_data_bus_0881_wide_signal ,
    output reg [31:0] \output_data_bus_0882_wide_signal ,
    output reg [31:0] \output_data_bus_0883_wide_signal ,
    output reg [31:0] \output_data_bus_0884_wide_signal ,
    output reg [31:0] \output_data_bus_0885_wide_signal ,
    output reg [31:0] \output_data_bus_0886_wide_signal ,
    output reg [31:0] \output_data_bus_0887_wide_signal ,
    output reg [31:0] \output_data_bus_0888_wide_signal ,
    output reg [31:0] \output_data_bus_0889_wide_signal ,
    output reg [31:0] \output_data_bus_0890_wide_signal ,
    output reg [31:0] \output_data_bus_0891_wide_signal ,
    output reg [31:0] \output_data_bus_0892_wide_signal ,
    output reg [31:0] \output_data_bus_0893_wide_signal ,
    output reg [31:0] \output_data_bus_0894_wide_signal ,
    output reg [31:0] \output_data_bus_0895_wide_signal ,
    output reg [31:0] \output_data_bus_0896_wide_signal ,
    output reg [31:0] \output_data_bus_0897_wide_signal ,
    output reg [31:0] \output_data_bus_0898_wide_signal ,
    output reg [31:0] \output_data_bus_0899_wide_signal ,
    output reg [31:0] \output_data_bus_0900_wide_signal ,
    output reg [31:0] \output_data_bus_0901_wide_signal ,
    output reg [31:0] \output_data_bus_0902_wide_signal ,
    output reg [31:0] \output_data_bus_0903_wide_signal ,
    output reg [31:0] \output_data_bus_0904_wide_signal ,
    output reg [31:0] \output_data_bus_0905_wide_signal ,
    output reg [31:0] \output_data_bus_0906_wide_signal ,
    output reg [31:0] \output_data_bus_0907_wide_signal ,
    output reg [31:0] \output_data_bus_0908_wide_signal ,
    output reg [31:0] \output_data_bus_0909_wide_signal ,
    output reg [31:0] \output_data_bus_0910_wide_signal ,
    output reg [31:0] \output_data_bus_0911_wide_signal ,
    output reg [31:0] \output_data_bus_0912_wide_signal ,
    output reg [31:0] \output_data_bus_0913_wide_signal ,
    output reg [31:0] \output_data_bus_0914_wide_signal ,
    output reg [31:0] \output_data_bus_0915_wide_signal ,
    output reg [31:0] \output_data_bus_0916_wide_signal ,
    output reg [31:0] \output_data_bus_0917_wide_signal ,
    output reg [31:0] \output_data_bus_0918_wide_signal ,
    output reg [31:0] \output_data_bus_0919_wide_signal ,
    output reg [31:0] \output_data_bus_0920_wide_signal ,
    output reg [31:0] \output_data_bus_0921_wide_signal ,
    output reg [31:0] \output_data_bus_0922_wide_signal ,
    output reg [31:0] \output_data_bus_0923_wide_signal ,
    output reg [31:0] \output_data_bus_0924_wide_signal ,
    output reg [31:0] \output_data_bus_0925_wide_signal ,
    output reg [31:0] \output_data_bus_0926_wide_signal ,
    output reg [31:0] \output_data_bus_0927_wide_signal ,
    output reg [31:0] \output_data_bus_0928_wide_signal ,
    output reg [31:0] \output_data_bus_0929_wide_signal ,
    output reg [31:0] \output_data_bus_0930_wide_signal ,
    output reg [31:0] \output_data_bus_0931_wide_signal ,
    output reg [31:0] \output_data_bus_0932_wide_signal ,
    output reg [31:0] \output_data_bus_0933_wide_signal ,
    output reg [31:0] \output_data_bus_0934_wide_signal ,
    output reg [31:0] \output_data_bus_0935_wide_signal ,
    output reg [31:0] \output_data_bus_0936_wide_signal ,
    output reg [31:0] \output_data_bus_0937_wide_signal ,
    output reg [31:0] \output_data_bus_0938_wide_signal ,
    output reg [31:0] \output_data_bus_0939_wide_signal ,
    output reg [31:0] \output_data_bus_0940_wide_signal ,
    output reg [31:0] \output_data_bus_0941_wide_signal ,
    output reg [31:0] \output_data_bus_0942_wide_signal ,
    output reg [31:0] \output_data_bus_0943_wide_signal ,
    output reg [31:0] \output_data_bus_0944_wide_signal ,
    output reg [31:0] \output_data_bus_0945_wide_signal ,
    output reg [31:0] \output_data_bus_0946_wide_signal ,
    output reg [31:0] \output_data_bus_0947_wide_signal ,
    output reg [31:0] \output_data_bus_0948_wide_signal ,
    output reg [31:0] \output_data_bus_0949_wide_signal ,
    output reg [31:0] \output_data_bus_0950_wide_signal ,
    output reg [31:0] \output_data_bus_0951_wide_signal ,
    output reg [31:0] \output_data_bus_0952_wide_signal ,
    output reg [31:0] \output_data_bus_0953_wide_signal ,
    output reg [31:0] \output_data_bus_0954_wide_signal ,
    output reg [31:0] \output_data_bus_0955_wide_signal ,
    output reg [31:0] \output_data_bus_0956_wide_signal ,
    output reg [31:0] \output_data_bus_0957_wide_signal ,
    output reg [31:0] \output_data_bus_0958_wide_signal ,
    output reg [31:0] \output_data_bus_0959_wide_signal ,
    output reg [31:0] \output_data_bus_0960_wide_signal ,
    output reg [31:0] \output_data_bus_0961_wide_signal ,
    output reg [31:0] \output_data_bus_0962_wide_signal ,
    output reg [31:0] \output_data_bus_0963_wide_signal ,
    output reg [31:0] \output_data_bus_0964_wide_signal ,
    output reg [31:0] \output_data_bus_0965_wide_signal ,
    output reg [31:0] \output_data_bus_0966_wide_signal ,
    output reg [31:0] \output_data_bus_0967_wide_signal ,
    output reg [31:0] \output_data_bus_0968_wide_signal ,
    output reg [31:0] \output_data_bus_0969_wide_signal ,
    output reg [31:0] \output_data_bus_0970_wide_signal ,
    output reg [31:0] \output_data_bus_0971_wide_signal ,
    output reg [31:0] \output_data_bus_0972_wide_signal ,
    output reg [31:0] \output_data_bus_0973_wide_signal ,
    output reg [31:0] \output_data_bus_0974_wide_signal ,
    output reg [31:0] \output_data_bus_0975_wide_signal ,
    output reg [31:0] \output_data_bus_0976_wide_signal ,
    output reg [31:0] \output_data_bus_0977_wide_signal ,
    output reg [31:0] \output_data_bus_0978_wide_signal ,
    output reg [31:0] \output_data_bus_0979_wide_signal ,
    output reg [31:0] \output_data_bus_0980_wide_signal ,
    output reg [31:0] \output_data_bus_0981_wide_signal ,
    output reg [31:0] \output_data_bus_0982_wide_signal ,
    output reg [31:0] \output_data_bus_0983_wide_signal ,
    output reg [31:0] \output_data_bus_0984_wide_signal ,
    output reg [31:0] \output_data_bus_0985_wide_signal ,
    output reg [31:0] \output_data_bus_0986_wide_signal ,
    output reg [31:0] \output_data_bus_0987_wide_signal ,
    output reg [31:0] \output_data_bus_0988_wide_signal ,
    output reg [31:0] \output_data_bus_0989_wide_signal ,
    output reg [31:0] \output_data_bus_0990_wide_signal ,
    output reg [31:0] \output_data_bus_0991_wide_signal ,
    output reg [31:0] \output_data_bus_0992_wide_signal ,
    output reg [31:0] \output_data_bus_0993_wide_signal ,
    output reg [31:0] \output_data_bus_0994_wide_signal ,
    output reg [31:0] \output_data_bus_0995_wide_signal ,
    output reg [31:0] \output_data_bus_0996_wide_signal ,
    output reg [31:0] \output_data_bus_0997_wide_signal ,
    output reg [31:0] \output_data_bus_0998_wide_signal ,
    output reg [31:0] \output_data_bus_0999_wide_signal ,
    inout [63:0] \bidir_data_bus_0000_ultra_wide ,
    inout [63:0] \bidir_data_bus_0001_ultra_wide ,
    inout [63:0] \bidir_data_bus_0002_ultra_wide ,
    inout [63:0] \bidir_data_bus_0003_ultra_wide ,
    inout [63:0] \bidir_data_bus_0004_ultra_wide ,
    inout [63:0] \bidir_data_bus_0005_ultra_wide ,
    inout [63:0] \bidir_data_bus_0006_ultra_wide ,
    inout [63:0] \bidir_data_bus_0007_ultra_wide ,
    inout [63:0] \bidir_data_bus_0008_ultra_wide ,
    inout [63:0] \bidir_data_bus_0009_ultra_wide ,
    inout [63:0] \bidir_data_bus_0010_ultra_wide ,
    inout [63:0] \bidir_data_bus_0011_ultra_wide ,
    inout [63:0] \bidir_data_bus_0012_ultra_wide ,
    inout [63:0] \bidir_data_bus_0013_ultra_wide ,
    inout [63:0] \bidir_data_bus_0014_ultra_wide ,
    inout [63:0] \bidir_data_bus_0015_ultra_wide ,
    inout [63:0] \bidir_data_bus_0016_ultra_wide ,
    inout [63:0] \bidir_data_bus_0017_ultra_wide ,
    inout [63:0] \bidir_data_bus_0018_ultra_wide ,
    inout [63:0] \bidir_data_bus_0019_ultra_wide ,
    inout [63:0] \bidir_data_bus_0020_ultra_wide ,
    inout [63:0] \bidir_data_bus_0021_ultra_wide ,
    inout [63:0] \bidir_data_bus_0022_ultra_wide ,
    inout [63:0] \bidir_data_bus_0023_ultra_wide ,
    inout [63:0] \bidir_data_bus_0024_ultra_wide ,
    inout [63:0] \bidir_data_bus_0025_ultra_wide ,
    inout [63:0] \bidir_data_bus_0026_ultra_wide ,
    inout [63:0] \bidir_data_bus_0027_ultra_wide ,
    inout [63:0] \bidir_data_bus_0028_ultra_wide ,
    inout [63:0] \bidir_data_bus_0029_ultra_wide ,
    inout [63:0] \bidir_data_bus_0030_ultra_wide ,
    inout [63:0] \bidir_data_bus_0031_ultra_wide ,
    inout [63:0] \bidir_data_bus_0032_ultra_wide ,
    inout [63:0] \bidir_data_bus_0033_ultra_wide ,
    inout [63:0] \bidir_data_bus_0034_ultra_wide ,
    inout [63:0] \bidir_data_bus_0035_ultra_wide ,
    inout [63:0] \bidir_data_bus_0036_ultra_wide ,
    inout [63:0] \bidir_data_bus_0037_ultra_wide ,
    inout [63:0] \bidir_data_bus_0038_ultra_wide ,
    inout [63:0] \bidir_data_bus_0039_ultra_wide ,
    inout [63:0] \bidir_data_bus_0040_ultra_wide ,
    inout [63:0] \bidir_data_bus_0041_ultra_wide ,
    inout [63:0] \bidir_data_bus_0042_ultra_wide ,
    inout [63:0] \bidir_data_bus_0043_ultra_wide ,
    inout [63:0] \bidir_data_bus_0044_ultra_wide ,
    inout [63:0] \bidir_data_bus_0045_ultra_wide ,
    inout [63:0] \bidir_data_bus_0046_ultra_wide ,
    inout [63:0] \bidir_data_bus_0047_ultra_wide ,
    inout [63:0] \bidir_data_bus_0048_ultra_wide ,
    inout [63:0] \bidir_data_bus_0049_ultra_wide ,
    inout [63:0] \bidir_data_bus_0050_ultra_wide ,
    inout [63:0] \bidir_data_bus_0051_ultra_wide ,
    inout [63:0] \bidir_data_bus_0052_ultra_wide ,
    inout [63:0] \bidir_data_bus_0053_ultra_wide ,
    inout [63:0] \bidir_data_bus_0054_ultra_wide ,
    inout [63:0] \bidir_data_bus_0055_ultra_wide ,
    inout [63:0] \bidir_data_bus_0056_ultra_wide ,
    inout [63:0] \bidir_data_bus_0057_ultra_wide ,
    inout [63:0] \bidir_data_bus_0058_ultra_wide ,
    inout [63:0] \bidir_data_bus_0059_ultra_wide ,
    inout [63:0] \bidir_data_bus_0060_ultra_wide ,
    inout [63:0] \bidir_data_bus_0061_ultra_wide ,
    inout [63:0] \bidir_data_bus_0062_ultra_wide ,
    inout [63:0] \bidir_data_bus_0063_ultra_wide ,
    inout [63:0] \bidir_data_bus_0064_ultra_wide ,
    inout [63:0] \bidir_data_bus_0065_ultra_wide ,
    inout [63:0] \bidir_data_bus_0066_ultra_wide ,
    inout [63:0] \bidir_data_bus_0067_ultra_wide ,
    inout [63:0] \bidir_data_bus_0068_ultra_wide ,
    inout [63:0] \bidir_data_bus_0069_ultra_wide ,
    inout [63:0] \bidir_data_bus_0070_ultra_wide ,
    inout [63:0] \bidir_data_bus_0071_ultra_wide ,
    inout [63:0] \bidir_data_bus_0072_ultra_wide ,
    inout [63:0] \bidir_data_bus_0073_ultra_wide ,
    inout [63:0] \bidir_data_bus_0074_ultra_wide ,
    inout [63:0] \bidir_data_bus_0075_ultra_wide ,
    inout [63:0] \bidir_data_bus_0076_ultra_wide ,
    inout [63:0] \bidir_data_bus_0077_ultra_wide ,
    inout [63:0] \bidir_data_bus_0078_ultra_wide ,
    inout [63:0] \bidir_data_bus_0079_ultra_wide ,
    inout [63:0] \bidir_data_bus_0080_ultra_wide ,
    inout [63:0] \bidir_data_bus_0081_ultra_wide ,
    inout [63:0] \bidir_data_bus_0082_ultra_wide ,
    inout [63:0] \bidir_data_bus_0083_ultra_wide ,
    inout [63:0] \bidir_data_bus_0084_ultra_wide ,
    inout [63:0] \bidir_data_bus_0085_ultra_wide ,
    inout [63:0] \bidir_data_bus_0086_ultra_wide ,
    inout [63:0] \bidir_data_bus_0087_ultra_wide ,
    inout [63:0] \bidir_data_bus_0088_ultra_wide ,
    inout [63:0] \bidir_data_bus_0089_ultra_wide ,
    inout [63:0] \bidir_data_bus_0090_ultra_wide ,
    inout [63:0] \bidir_data_bus_0091_ultra_wide ,
    inout [63:0] \bidir_data_bus_0092_ultra_wide ,
    inout [63:0] \bidir_data_bus_0093_ultra_wide ,
    inout [63:0] \bidir_data_bus_0094_ultra_wide ,
    inout [63:0] \bidir_data_bus_0095_ultra_wide ,
    inout [63:0] \bidir_data_bus_0096_ultra_wide ,
    inout [63:0] \bidir_data_bus_0097_ultra_wide ,
    inout [63:0] \bidir_data_bus_0098_ultra_wide ,
    inout [63:0] \bidir_data_bus_0099_ultra_wide ,
    inout [63:0] \bidir_data_bus_0100_ultra_wide ,
    inout [63:0] \bidir_data_bus_0101_ultra_wide ,
    inout [63:0] \bidir_data_bus_0102_ultra_wide ,
    inout [63:0] \bidir_data_bus_0103_ultra_wide ,
    inout [63:0] \bidir_data_bus_0104_ultra_wide ,
    inout [63:0] \bidir_data_bus_0105_ultra_wide ,
    inout [63:0] \bidir_data_bus_0106_ultra_wide ,
    inout [63:0] \bidir_data_bus_0107_ultra_wide ,
    inout [63:0] \bidir_data_bus_0108_ultra_wide ,
    inout [63:0] \bidir_data_bus_0109_ultra_wide ,
    inout [63:0] \bidir_data_bus_0110_ultra_wide ,
    inout [63:0] \bidir_data_bus_0111_ultra_wide ,
    inout [63:0] \bidir_data_bus_0112_ultra_wide ,
    inout [63:0] \bidir_data_bus_0113_ultra_wide ,
    inout [63:0] \bidir_data_bus_0114_ultra_wide ,
    inout [63:0] \bidir_data_bus_0115_ultra_wide ,
    inout [63:0] \bidir_data_bus_0116_ultra_wide ,
    inout [63:0] \bidir_data_bus_0117_ultra_wide ,
    inout [63:0] \bidir_data_bus_0118_ultra_wide ,
    inout [63:0] \bidir_data_bus_0119_ultra_wide ,
    inout [63:0] \bidir_data_bus_0120_ultra_wide ,
    inout [63:0] \bidir_data_bus_0121_ultra_wide ,
    inout [63:0] \bidir_data_bus_0122_ultra_wide ,
    inout [63:0] \bidir_data_bus_0123_ultra_wide ,
    inout [63:0] \bidir_data_bus_0124_ultra_wide ,
    inout [63:0] \bidir_data_bus_0125_ultra_wide ,
    inout [63:0] \bidir_data_bus_0126_ultra_wide ,
    inout [63:0] \bidir_data_bus_0127_ultra_wide ,
    inout [63:0] \bidir_data_bus_0128_ultra_wide ,
    inout [63:0] \bidir_data_bus_0129_ultra_wide ,
    inout [63:0] \bidir_data_bus_0130_ultra_wide ,
    inout [63:0] \bidir_data_bus_0131_ultra_wide ,
    inout [63:0] \bidir_data_bus_0132_ultra_wide ,
    inout [63:0] \bidir_data_bus_0133_ultra_wide ,
    inout [63:0] \bidir_data_bus_0134_ultra_wide ,
    inout [63:0] \bidir_data_bus_0135_ultra_wide ,
    inout [63:0] \bidir_data_bus_0136_ultra_wide ,
    inout [63:0] \bidir_data_bus_0137_ultra_wide ,
    inout [63:0] \bidir_data_bus_0138_ultra_wide ,
    inout [63:0] \bidir_data_bus_0139_ultra_wide ,
    inout [63:0] \bidir_data_bus_0140_ultra_wide ,
    inout [63:0] \bidir_data_bus_0141_ultra_wide ,
    inout [63:0] \bidir_data_bus_0142_ultra_wide ,
    inout [63:0] \bidir_data_bus_0143_ultra_wide ,
    inout [63:0] \bidir_data_bus_0144_ultra_wide ,
    inout [63:0] \bidir_data_bus_0145_ultra_wide ,
    inout [63:0] \bidir_data_bus_0146_ultra_wide ,
    inout [63:0] \bidir_data_bus_0147_ultra_wide ,
    inout [63:0] \bidir_data_bus_0148_ultra_wide ,
    inout [63:0] \bidir_data_bus_0149_ultra_wide ,
    inout [63:0] \bidir_data_bus_0150_ultra_wide ,
    inout [63:0] \bidir_data_bus_0151_ultra_wide ,
    inout [63:0] \bidir_data_bus_0152_ultra_wide ,
    inout [63:0] \bidir_data_bus_0153_ultra_wide ,
    inout [63:0] \bidir_data_bus_0154_ultra_wide ,
    inout [63:0] \bidir_data_bus_0155_ultra_wide ,
    inout [63:0] \bidir_data_bus_0156_ultra_wide ,
    inout [63:0] \bidir_data_bus_0157_ultra_wide ,
    inout [63:0] \bidir_data_bus_0158_ultra_wide ,
    inout [63:0] \bidir_data_bus_0159_ultra_wide ,
    inout [63:0] \bidir_data_bus_0160_ultra_wide ,
    inout [63:0] \bidir_data_bus_0161_ultra_wide ,
    inout [63:0] \bidir_data_bus_0162_ultra_wide ,
    inout [63:0] \bidir_data_bus_0163_ultra_wide ,
    inout [63:0] \bidir_data_bus_0164_ultra_wide ,
    inout [63:0] \bidir_data_bus_0165_ultra_wide ,
    inout [63:0] \bidir_data_bus_0166_ultra_wide ,
    inout [63:0] \bidir_data_bus_0167_ultra_wide ,
    inout [63:0] \bidir_data_bus_0168_ultra_wide ,
    inout [63:0] \bidir_data_bus_0169_ultra_wide ,
    inout [63:0] \bidir_data_bus_0170_ultra_wide ,
    inout [63:0] \bidir_data_bus_0171_ultra_wide ,
    inout [63:0] \bidir_data_bus_0172_ultra_wide ,
    inout [63:0] \bidir_data_bus_0173_ultra_wide ,
    inout [63:0] \bidir_data_bus_0174_ultra_wide ,
    inout [63:0] \bidir_data_bus_0175_ultra_wide ,
    inout [63:0] \bidir_data_bus_0176_ultra_wide ,
    inout [63:0] \bidir_data_bus_0177_ultra_wide ,
    inout [63:0] \bidir_data_bus_0178_ultra_wide ,
    inout [63:0] \bidir_data_bus_0179_ultra_wide ,
    inout [63:0] \bidir_data_bus_0180_ultra_wide ,
    inout [63:0] \bidir_data_bus_0181_ultra_wide ,
    inout [63:0] \bidir_data_bus_0182_ultra_wide ,
    inout [63:0] \bidir_data_bus_0183_ultra_wide ,
    inout [63:0] \bidir_data_bus_0184_ultra_wide ,
    inout [63:0] \bidir_data_bus_0185_ultra_wide ,
    inout [63:0] \bidir_data_bus_0186_ultra_wide ,
    inout [63:0] \bidir_data_bus_0187_ultra_wide ,
    inout [63:0] \bidir_data_bus_0188_ultra_wide ,
    inout [63:0] \bidir_data_bus_0189_ultra_wide ,
    inout [63:0] \bidir_data_bus_0190_ultra_wide ,
    inout [63:0] \bidir_data_bus_0191_ultra_wide ,
    inout [63:0] \bidir_data_bus_0192_ultra_wide ,
    inout [63:0] \bidir_data_bus_0193_ultra_wide ,
    inout [63:0] \bidir_data_bus_0194_ultra_wide ,
    inout [63:0] \bidir_data_bus_0195_ultra_wide ,
    inout [63:0] \bidir_data_bus_0196_ultra_wide ,
    inout [63:0] \bidir_data_bus_0197_ultra_wide ,
    inout [63:0] \bidir_data_bus_0198_ultra_wide ,
    inout [63:0] \bidir_data_bus_0199_ultra_wide ,
    inout [63:0] \bidir_data_bus_0200_ultra_wide ,
    inout [63:0] \bidir_data_bus_0201_ultra_wide ,
    inout [63:0] \bidir_data_bus_0202_ultra_wide ,
    inout [63:0] \bidir_data_bus_0203_ultra_wide ,
    inout [63:0] \bidir_data_bus_0204_ultra_wide ,
    inout [63:0] \bidir_data_bus_0205_ultra_wide ,
    inout [63:0] \bidir_data_bus_0206_ultra_wide ,
    inout [63:0] \bidir_data_bus_0207_ultra_wide ,
    inout [63:0] \bidir_data_bus_0208_ultra_wide ,
    inout [63:0] \bidir_data_bus_0209_ultra_wide ,
    inout [63:0] \bidir_data_bus_0210_ultra_wide ,
    inout [63:0] \bidir_data_bus_0211_ultra_wide ,
    inout [63:0] \bidir_data_bus_0212_ultra_wide ,
    inout [63:0] \bidir_data_bus_0213_ultra_wide ,
    inout [63:0] \bidir_data_bus_0214_ultra_wide ,
    inout [63:0] \bidir_data_bus_0215_ultra_wide ,
    inout [63:0] \bidir_data_bus_0216_ultra_wide ,
    inout [63:0] \bidir_data_bus_0217_ultra_wide ,
    inout [63:0] \bidir_data_bus_0218_ultra_wide ,
    inout [63:0] \bidir_data_bus_0219_ultra_wide ,
    inout [63:0] \bidir_data_bus_0220_ultra_wide ,
    inout [63:0] \bidir_data_bus_0221_ultra_wide ,
    inout [63:0] \bidir_data_bus_0222_ultra_wide ,
    inout [63:0] \bidir_data_bus_0223_ultra_wide ,
    inout [63:0] \bidir_data_bus_0224_ultra_wide ,
    inout [63:0] \bidir_data_bus_0225_ultra_wide ,
    inout [63:0] \bidir_data_bus_0226_ultra_wide ,
    inout [63:0] \bidir_data_bus_0227_ultra_wide ,
    inout [63:0] \bidir_data_bus_0228_ultra_wide ,
    inout [63:0] \bidir_data_bus_0229_ultra_wide ,
    inout [63:0] \bidir_data_bus_0230_ultra_wide ,
    inout [63:0] \bidir_data_bus_0231_ultra_wide ,
    inout [63:0] \bidir_data_bus_0232_ultra_wide ,
    inout [63:0] \bidir_data_bus_0233_ultra_wide ,
    inout [63:0] \bidir_data_bus_0234_ultra_wide ,
    inout [63:0] \bidir_data_bus_0235_ultra_wide ,
    inout [63:0] \bidir_data_bus_0236_ultra_wide ,
    inout [63:0] \bidir_data_bus_0237_ultra_wide ,
    inout [63:0] \bidir_data_bus_0238_ultra_wide ,
    inout [63:0] \bidir_data_bus_0239_ultra_wide ,
    inout [63:0] \bidir_data_bus_0240_ultra_wide ,
    inout [63:0] \bidir_data_bus_0241_ultra_wide ,
    inout [63:0] \bidir_data_bus_0242_ultra_wide ,
    inout [63:0] \bidir_data_bus_0243_ultra_wide ,
    inout [63:0] \bidir_data_bus_0244_ultra_wide ,
    inout [63:0] \bidir_data_bus_0245_ultra_wide ,
    inout [63:0] \bidir_data_bus_0246_ultra_wide ,
    inout [63:0] \bidir_data_bus_0247_ultra_wide ,
    inout [63:0] \bidir_data_bus_0248_ultra_wide ,
    inout [63:0] \bidir_data_bus_0249_ultra_wide ,
    inout [63:0] \bidir_data_bus_0250_ultra_wide ,
    inout [63:0] \bidir_data_bus_0251_ultra_wide ,
    inout [63:0] \bidir_data_bus_0252_ultra_wide ,
    inout [63:0] \bidir_data_bus_0253_ultra_wide ,
    inout [63:0] \bidir_data_bus_0254_ultra_wide ,
    inout [63:0] \bidir_data_bus_0255_ultra_wide ,
    inout [63:0] \bidir_data_bus_0256_ultra_wide ,
    inout [63:0] \bidir_data_bus_0257_ultra_wide ,
    inout [63:0] \bidir_data_bus_0258_ultra_wide ,
    inout [63:0] \bidir_data_bus_0259_ultra_wide ,
    inout [63:0] \bidir_data_bus_0260_ultra_wide ,
    inout [63:0] \bidir_data_bus_0261_ultra_wide ,
    inout [63:0] \bidir_data_bus_0262_ultra_wide ,
    inout [63:0] \bidir_data_bus_0263_ultra_wide ,
    inout [63:0] \bidir_data_bus_0264_ultra_wide ,
    inout [63:0] \bidir_data_bus_0265_ultra_wide ,
    inout [63:0] \bidir_data_bus_0266_ultra_wide ,
    inout [63:0] \bidir_data_bus_0267_ultra_wide ,
    inout [63:0] \bidir_data_bus_0268_ultra_wide ,
    inout [63:0] \bidir_data_bus_0269_ultra_wide ,
    inout [63:0] \bidir_data_bus_0270_ultra_wide ,
    inout [63:0] \bidir_data_bus_0271_ultra_wide ,
    inout [63:0] \bidir_data_bus_0272_ultra_wide ,
    inout [63:0] \bidir_data_bus_0273_ultra_wide ,
    inout [63:0] \bidir_data_bus_0274_ultra_wide ,
    inout [63:0] \bidir_data_bus_0275_ultra_wide ,
    inout [63:0] \bidir_data_bus_0276_ultra_wide ,
    inout [63:0] \bidir_data_bus_0277_ultra_wide ,
    inout [63:0] \bidir_data_bus_0278_ultra_wide ,
    inout [63:0] \bidir_data_bus_0279_ultra_wide ,
    inout [63:0] \bidir_data_bus_0280_ultra_wide ,
    inout [63:0] \bidir_data_bus_0281_ultra_wide ,
    inout [63:0] \bidir_data_bus_0282_ultra_wide ,
    inout [63:0] \bidir_data_bus_0283_ultra_wide ,
    inout [63:0] \bidir_data_bus_0284_ultra_wide ,
    inout [63:0] \bidir_data_bus_0285_ultra_wide ,
    inout [63:0] \bidir_data_bus_0286_ultra_wide ,
    inout [63:0] \bidir_data_bus_0287_ultra_wide ,
    inout [63:0] \bidir_data_bus_0288_ultra_wide ,
    inout [63:0] \bidir_data_bus_0289_ultra_wide ,
    inout [63:0] \bidir_data_bus_0290_ultra_wide ,
    inout [63:0] \bidir_data_bus_0291_ultra_wide ,
    inout [63:0] \bidir_data_bus_0292_ultra_wide ,
    inout [63:0] \bidir_data_bus_0293_ultra_wide ,
    inout [63:0] \bidir_data_bus_0294_ultra_wide ,
    inout [63:0] \bidir_data_bus_0295_ultra_wide ,
    inout [63:0] \bidir_data_bus_0296_ultra_wide ,
    inout [63:0] \bidir_data_bus_0297_ultra_wide ,
    inout [63:0] \bidir_data_bus_0298_ultra_wide ,
    inout [63:0] \bidir_data_bus_0299_ultra_wide ,
    inout [63:0] \bidir_data_bus_0300_ultra_wide ,
    inout [63:0] \bidir_data_bus_0301_ultra_wide ,
    inout [63:0] \bidir_data_bus_0302_ultra_wide ,
    inout [63:0] \bidir_data_bus_0303_ultra_wide ,
    inout [63:0] \bidir_data_bus_0304_ultra_wide ,
    inout [63:0] \bidir_data_bus_0305_ultra_wide ,
    inout [63:0] \bidir_data_bus_0306_ultra_wide ,
    inout [63:0] \bidir_data_bus_0307_ultra_wide ,
    inout [63:0] \bidir_data_bus_0308_ultra_wide ,
    inout [63:0] \bidir_data_bus_0309_ultra_wide ,
    inout [63:0] \bidir_data_bus_0310_ultra_wide ,
    inout [63:0] \bidir_data_bus_0311_ultra_wide ,
    inout [63:0] \bidir_data_bus_0312_ultra_wide ,
    inout [63:0] \bidir_data_bus_0313_ultra_wide ,
    inout [63:0] \bidir_data_bus_0314_ultra_wide ,
    inout [63:0] \bidir_data_bus_0315_ultra_wide ,
    inout [63:0] \bidir_data_bus_0316_ultra_wide ,
    inout [63:0] \bidir_data_bus_0317_ultra_wide ,
    inout [63:0] \bidir_data_bus_0318_ultra_wide ,
    inout [63:0] \bidir_data_bus_0319_ultra_wide ,
    inout [63:0] \bidir_data_bus_0320_ultra_wide ,
    inout [63:0] \bidir_data_bus_0321_ultra_wide ,
    inout [63:0] \bidir_data_bus_0322_ultra_wide ,
    inout [63:0] \bidir_data_bus_0323_ultra_wide ,
    inout [63:0] \bidir_data_bus_0324_ultra_wide ,
    inout [63:0] \bidir_data_bus_0325_ultra_wide ,
    inout [63:0] \bidir_data_bus_0326_ultra_wide ,
    inout [63:0] \bidir_data_bus_0327_ultra_wide ,
    inout [63:0] \bidir_data_bus_0328_ultra_wide ,
    inout [63:0] \bidir_data_bus_0329_ultra_wide ,
    inout [63:0] \bidir_data_bus_0330_ultra_wide ,
    inout [63:0] \bidir_data_bus_0331_ultra_wide ,
    inout [63:0] \bidir_data_bus_0332_ultra_wide ,
    inout [63:0] \bidir_data_bus_0333_ultra_wide ,
    inout [63:0] \bidir_data_bus_0334_ultra_wide ,
    inout [63:0] \bidir_data_bus_0335_ultra_wide ,
    inout [63:0] \bidir_data_bus_0336_ultra_wide ,
    inout [63:0] \bidir_data_bus_0337_ultra_wide ,
    inout [63:0] \bidir_data_bus_0338_ultra_wide ,
    inout [63:0] \bidir_data_bus_0339_ultra_wide ,
    inout [63:0] \bidir_data_bus_0340_ultra_wide ,
    inout [63:0] \bidir_data_bus_0341_ultra_wide ,
    inout [63:0] \bidir_data_bus_0342_ultra_wide ,
    inout [63:0] \bidir_data_bus_0343_ultra_wide ,
    inout [63:0] \bidir_data_bus_0344_ultra_wide ,
    inout [63:0] \bidir_data_bus_0345_ultra_wide ,
    inout [63:0] \bidir_data_bus_0346_ultra_wide ,
    inout [63:0] \bidir_data_bus_0347_ultra_wide ,
    inout [63:0] \bidir_data_bus_0348_ultra_wide ,
    inout [63:0] \bidir_data_bus_0349_ultra_wide ,
    inout [63:0] \bidir_data_bus_0350_ultra_wide ,
    inout [63:0] \bidir_data_bus_0351_ultra_wide ,
    inout [63:0] \bidir_data_bus_0352_ultra_wide ,
    inout [63:0] \bidir_data_bus_0353_ultra_wide ,
    inout [63:0] \bidir_data_bus_0354_ultra_wide ,
    inout [63:0] \bidir_data_bus_0355_ultra_wide ,
    inout [63:0] \bidir_data_bus_0356_ultra_wide ,
    inout [63:0] \bidir_data_bus_0357_ultra_wide ,
    inout [63:0] \bidir_data_bus_0358_ultra_wide ,
    inout [63:0] \bidir_data_bus_0359_ultra_wide ,
    inout [63:0] \bidir_data_bus_0360_ultra_wide ,
    inout [63:0] \bidir_data_bus_0361_ultra_wide ,
    inout [63:0] \bidir_data_bus_0362_ultra_wide ,
    inout [63:0] \bidir_data_bus_0363_ultra_wide ,
    inout [63:0] \bidir_data_bus_0364_ultra_wide ,
    inout [63:0] \bidir_data_bus_0365_ultra_wide ,
    inout [63:0] \bidir_data_bus_0366_ultra_wide ,
    inout [63:0] \bidir_data_bus_0367_ultra_wide ,
    inout [63:0] \bidir_data_bus_0368_ultra_wide ,
    inout [63:0] \bidir_data_bus_0369_ultra_wide ,
    inout [63:0] \bidir_data_bus_0370_ultra_wide ,
    inout [63:0] \bidir_data_bus_0371_ultra_wide ,
    inout [63:0] \bidir_data_bus_0372_ultra_wide ,
    inout [63:0] \bidir_data_bus_0373_ultra_wide ,
    inout [63:0] \bidir_data_bus_0374_ultra_wide ,
    inout [63:0] \bidir_data_bus_0375_ultra_wide ,
    inout [63:0] \bidir_data_bus_0376_ultra_wide ,
    inout [63:0] \bidir_data_bus_0377_ultra_wide ,
    inout [63:0] \bidir_data_bus_0378_ultra_wide ,
    inout [63:0] \bidir_data_bus_0379_ultra_wide ,
    inout [63:0] \bidir_data_bus_0380_ultra_wide ,
    inout [63:0] \bidir_data_bus_0381_ultra_wide ,
    inout [63:0] \bidir_data_bus_0382_ultra_wide ,
    inout [63:0] \bidir_data_bus_0383_ultra_wide ,
    inout [63:0] \bidir_data_bus_0384_ultra_wide ,
    inout [63:0] \bidir_data_bus_0385_ultra_wide ,
    inout [63:0] \bidir_data_bus_0386_ultra_wide ,
    inout [63:0] \bidir_data_bus_0387_ultra_wide ,
    inout [63:0] \bidir_data_bus_0388_ultra_wide ,
    inout [63:0] \bidir_data_bus_0389_ultra_wide ,
    inout [63:0] \bidir_data_bus_0390_ultra_wide ,
    inout [63:0] \bidir_data_bus_0391_ultra_wide ,
    inout [63:0] \bidir_data_bus_0392_ultra_wide ,
    inout [63:0] \bidir_data_bus_0393_ultra_wide ,
    inout [63:0] \bidir_data_bus_0394_ultra_wide ,
    inout [63:0] \bidir_data_bus_0395_ultra_wide ,
    inout [63:0] \bidir_data_bus_0396_ultra_wide ,
    inout [63:0] \bidir_data_bus_0397_ultra_wide ,
    inout [63:0] \bidir_data_bus_0398_ultra_wide ,
    inout [63:0] \bidir_data_bus_0399_ultra_wide ,
    inout [63:0] \bidir_data_bus_0400_ultra_wide ,
    inout [63:0] \bidir_data_bus_0401_ultra_wide ,
    inout [63:0] \bidir_data_bus_0402_ultra_wide ,
    inout [63:0] \bidir_data_bus_0403_ultra_wide ,
    inout [63:0] \bidir_data_bus_0404_ultra_wide ,
    inout [63:0] \bidir_data_bus_0405_ultra_wide ,
    inout [63:0] \bidir_data_bus_0406_ultra_wide ,
    inout [63:0] \bidir_data_bus_0407_ultra_wide ,
    inout [63:0] \bidir_data_bus_0408_ultra_wide ,
    inout [63:0] \bidir_data_bus_0409_ultra_wide ,
    inout [63:0] \bidir_data_bus_0410_ultra_wide ,
    inout [63:0] \bidir_data_bus_0411_ultra_wide ,
    inout [63:0] \bidir_data_bus_0412_ultra_wide ,
    inout [63:0] \bidir_data_bus_0413_ultra_wide ,
    inout [63:0] \bidir_data_bus_0414_ultra_wide ,
    inout [63:0] \bidir_data_bus_0415_ultra_wide ,
    inout [63:0] \bidir_data_bus_0416_ultra_wide ,
    inout [63:0] \bidir_data_bus_0417_ultra_wide ,
    inout [63:0] \bidir_data_bus_0418_ultra_wide ,
    inout [63:0] \bidir_data_bus_0419_ultra_wide ,
    inout [63:0] \bidir_data_bus_0420_ultra_wide ,
    inout [63:0] \bidir_data_bus_0421_ultra_wide ,
    inout [63:0] \bidir_data_bus_0422_ultra_wide ,
    inout [63:0] \bidir_data_bus_0423_ultra_wide ,
    inout [63:0] \bidir_data_bus_0424_ultra_wide ,
    inout [63:0] \bidir_data_bus_0425_ultra_wide ,
    inout [63:0] \bidir_data_bus_0426_ultra_wide ,
    inout [63:0] \bidir_data_bus_0427_ultra_wide ,
    inout [63:0] \bidir_data_bus_0428_ultra_wide ,
    inout [63:0] \bidir_data_bus_0429_ultra_wide ,
    inout [63:0] \bidir_data_bus_0430_ultra_wide ,
    inout [63:0] \bidir_data_bus_0431_ultra_wide ,
    inout [63:0] \bidir_data_bus_0432_ultra_wide ,
    inout [63:0] \bidir_data_bus_0433_ultra_wide ,
    inout [63:0] \bidir_data_bus_0434_ultra_wide ,
    inout [63:0] \bidir_data_bus_0435_ultra_wide ,
    inout [63:0] \bidir_data_bus_0436_ultra_wide ,
    inout [63:0] \bidir_data_bus_0437_ultra_wide ,
    inout [63:0] \bidir_data_bus_0438_ultra_wide ,
    inout [63:0] \bidir_data_bus_0439_ultra_wide ,
    inout [63:0] \bidir_data_bus_0440_ultra_wide ,
    inout [63:0] \bidir_data_bus_0441_ultra_wide ,
    inout [63:0] \bidir_data_bus_0442_ultra_wide ,
    inout [63:0] \bidir_data_bus_0443_ultra_wide ,
    inout [63:0] \bidir_data_bus_0444_ultra_wide ,
    inout [63:0] \bidir_data_bus_0445_ultra_wide ,
    inout [63:0] \bidir_data_bus_0446_ultra_wide ,
    inout [63:0] \bidir_data_bus_0447_ultra_wide ,
    inout [63:0] \bidir_data_bus_0448_ultra_wide ,
    inout [63:0] \bidir_data_bus_0449_ultra_wide ,
    inout [63:0] \bidir_data_bus_0450_ultra_wide ,
    inout [63:0] \bidir_data_bus_0451_ultra_wide ,
    inout [63:0] \bidir_data_bus_0452_ultra_wide ,
    inout [63:0] \bidir_data_bus_0453_ultra_wide ,
    inout [63:0] \bidir_data_bus_0454_ultra_wide ,
    inout [63:0] \bidir_data_bus_0455_ultra_wide ,
    inout [63:0] \bidir_data_bus_0456_ultra_wide ,
    inout [63:0] \bidir_data_bus_0457_ultra_wide ,
    inout [63:0] \bidir_data_bus_0458_ultra_wide ,
    inout [63:0] \bidir_data_bus_0459_ultra_wide ,
    inout [63:0] \bidir_data_bus_0460_ultra_wide ,
    inout [63:0] \bidir_data_bus_0461_ultra_wide ,
    inout [63:0] \bidir_data_bus_0462_ultra_wide ,
    inout [63:0] \bidir_data_bus_0463_ultra_wide ,
    inout [63:0] \bidir_data_bus_0464_ultra_wide ,
    inout [63:0] \bidir_data_bus_0465_ultra_wide ,
    inout [63:0] \bidir_data_bus_0466_ultra_wide ,
    inout [63:0] \bidir_data_bus_0467_ultra_wide ,
    inout [63:0] \bidir_data_bus_0468_ultra_wide ,
    inout [63:0] \bidir_data_bus_0469_ultra_wide ,
    inout [63:0] \bidir_data_bus_0470_ultra_wide ,
    inout [63:0] \bidir_data_bus_0471_ultra_wide ,
    inout [63:0] \bidir_data_bus_0472_ultra_wide ,
    inout [63:0] \bidir_data_bus_0473_ultra_wide ,
    inout [63:0] \bidir_data_bus_0474_ultra_wide ,
    inout [63:0] \bidir_data_bus_0475_ultra_wide ,
    inout [63:0] \bidir_data_bus_0476_ultra_wide ,
    inout [63:0] \bidir_data_bus_0477_ultra_wide ,
    inout [63:0] \bidir_data_bus_0478_ultra_wide ,
    inout [63:0] \bidir_data_bus_0479_ultra_wide ,
    inout [63:0] \bidir_data_bus_0480_ultra_wide ,
    inout [63:0] \bidir_data_bus_0481_ultra_wide ,
    inout [63:0] \bidir_data_bus_0482_ultra_wide ,
    inout [63:0] \bidir_data_bus_0483_ultra_wide ,
    inout [63:0] \bidir_data_bus_0484_ultra_wide ,
    inout [63:0] \bidir_data_bus_0485_ultra_wide ,
    inout [63:0] \bidir_data_bus_0486_ultra_wide ,
    inout [63:0] \bidir_data_bus_0487_ultra_wide ,
    inout [63:0] \bidir_data_bus_0488_ultra_wide ,
    inout [63:0] \bidir_data_bus_0489_ultra_wide ,
    inout [63:0] \bidir_data_bus_0490_ultra_wide ,
    inout [63:0] \bidir_data_bus_0491_ultra_wide ,
    inout [63:0] \bidir_data_bus_0492_ultra_wide ,
    inout [63:0] \bidir_data_bus_0493_ultra_wide ,
    inout [63:0] \bidir_data_bus_0494_ultra_wide ,
    inout [63:0] \bidir_data_bus_0495_ultra_wide ,
    inout [63:0] \bidir_data_bus_0496_ultra_wide ,
    inout [63:0] \bidir_data_bus_0497_ultra_wide ,
    inout [63:0] \bidir_data_bus_0498_ultra_wide ,
    inout [63:0] \bidir_data_bus_0499_ultra_wide 
);

// Internal registers for complex logic
reg [127:0] \internal_reg_bank_000_storage ;
reg [127:0] \internal_reg_bank_001_storage ;
reg [127:0] \internal_reg_bank_002_storage ;
reg [127:0] \internal_reg_bank_003_storage ;
reg [127:0] \internal_reg_bank_004_storage ;
reg [127:0] \internal_reg_bank_005_storage ;
reg [127:0] \internal_reg_bank_006_storage ;
reg [127:0] \internal_reg_bank_007_storage ;
reg [127:0] \internal_reg_bank_008_storage ;
reg [127:0] \internal_reg_bank_009_storage ;
reg [127:0] \internal_reg_bank_010_storage ;
reg [127:0] \internal_reg_bank_011_storage ;
reg [127:0] \internal_reg_bank_012_storage ;
reg [127:0] \internal_reg_bank_013_storage ;
reg [127:0] \internal_reg_bank_014_storage ;
reg [127:0] \internal_reg_bank_015_storage ;
reg [127:0] \internal_reg_bank_016_storage ;
reg [127:0] \internal_reg_bank_017_storage ;
reg [127:0] \internal_reg_bank_018_storage ;
reg [127:0] \internal_reg_bank_019_storage ;
reg [127:0] \internal_reg_bank_020_storage ;
reg [127:0] \internal_reg_bank_021_storage ;
reg [127:0] \internal_reg_bank_022_storage ;
reg [127:0] \internal_reg_bank_023_storage ;
reg [127:0] \internal_reg_bank_024_storage ;
reg [127:0] \internal_reg_bank_025_storage ;
reg [127:0] \internal_reg_bank_026_storage ;
reg [127:0] \internal_reg_bank_027_storage ;
reg [127:0] \internal_reg_bank_028_storage ;
reg [127:0] \internal_reg_bank_029_storage ;
reg [127:0] \internal_reg_bank_030_storage ;
reg [127:0] \internal_reg_bank_031_storage ;
reg [127:0] \internal_reg_bank_032_storage ;
reg [127:0] \internal_reg_bank_033_storage ;
reg [127:0] \internal_reg_bank_034_storage ;
reg [127:0] \internal_reg_bank_035_storage ;
reg [127:0] \internal_reg_bank_036_storage ;
reg [127:0] \internal_reg_bank_037_storage ;
reg [127:0] \internal_reg_bank_038_storage ;
reg [127:0] \internal_reg_bank_039_storage ;
reg [127:0] \internal_reg_bank_040_storage ;
reg [127:0] \internal_reg_bank_041_storage ;
reg [127:0] \internal_reg_bank_042_storage ;
reg [127:0] \internal_reg_bank_043_storage ;
reg [127:0] \internal_reg_bank_044_storage ;
reg [127:0] \internal_reg_bank_045_storage ;
reg [127:0] \internal_reg_bank_046_storage ;
reg [127:0] \internal_reg_bank_047_storage ;
reg [127:0] \internal_reg_bank_048_storage ;
reg [127:0] \internal_reg_bank_049_storage ;
reg [127:0] \internal_reg_bank_050_storage ;
reg [127:0] \internal_reg_bank_051_storage ;
reg [127:0] \internal_reg_bank_052_storage ;
reg [127:0] \internal_reg_bank_053_storage ;
reg [127:0] \internal_reg_bank_054_storage ;
reg [127:0] \internal_reg_bank_055_storage ;
reg [127:0] \internal_reg_bank_056_storage ;
reg [127:0] \internal_reg_bank_057_storage ;
reg [127:0] \internal_reg_bank_058_storage ;
reg [127:0] \internal_reg_bank_059_storage ;
reg [127:0] \internal_reg_bank_060_storage ;
reg [127:0] \internal_reg_bank_061_storage ;
reg [127:0] \internal_reg_bank_062_storage ;
reg [127:0] \internal_reg_bank_063_storage ;
reg [127:0] \internal_reg_bank_064_storage ;
reg [127:0] \internal_reg_bank_065_storage ;
reg [127:0] \internal_reg_bank_066_storage ;
reg [127:0] \internal_reg_bank_067_storage ;
reg [127:0] \internal_reg_bank_068_storage ;
reg [127:0] \internal_reg_bank_069_storage ;
reg [127:0] \internal_reg_bank_070_storage ;
reg [127:0] \internal_reg_bank_071_storage ;
reg [127:0] \internal_reg_bank_072_storage ;
reg [127:0] \internal_reg_bank_073_storage ;
reg [127:0] \internal_reg_bank_074_storage ;
reg [127:0] \internal_reg_bank_075_storage ;
reg [127:0] \internal_reg_bank_076_storage ;
reg [127:0] \internal_reg_bank_077_storage ;
reg [127:0] \internal_reg_bank_078_storage ;
reg [127:0] \internal_reg_bank_079_storage ;
reg [127:0] \internal_reg_bank_080_storage ;
reg [127:0] \internal_reg_bank_081_storage ;
reg [127:0] \internal_reg_bank_082_storage ;
reg [127:0] \internal_reg_bank_083_storage ;
reg [127:0] \internal_reg_bank_084_storage ;
reg [127:0] \internal_reg_bank_085_storage ;
reg [127:0] \internal_reg_bank_086_storage ;
reg [127:0] \internal_reg_bank_087_storage ;
reg [127:0] \internal_reg_bank_088_storage ;
reg [127:0] \internal_reg_bank_089_storage ;
reg [127:0] \internal_reg_bank_090_storage ;
reg [127:0] \internal_reg_bank_091_storage ;
reg [127:0] \internal_reg_bank_092_storage ;
reg [127:0] \internal_reg_bank_093_storage ;
reg [127:0] \internal_reg_bank_094_storage ;
reg [127:0] \internal_reg_bank_095_storage ;
reg [127:0] \internal_reg_bank_096_storage ;
reg [127:0] \internal_reg_bank_097_storage ;
reg [127:0] \internal_reg_bank_098_storage ;
reg [127:0] \internal_reg_bank_099_storage ;

// Deep nested generate blocks
genvar i, j, k;
generate
    for (i = 0; i < 32; i = i + 1) begin : gen_level_1
        for (j = 0; j < 16; j = j + 1) begin : gen_level_2
            for (k = 0; k < 8; k = k + 1) begin : gen_level_3
                reg [15:0] \nested_reg_array ;
            end
        end
    end
endgenerate

// Complex always block with many signals
always @(posedge clk_main_200mhz or negedge reset_n) begin
    if (!reset_n) begin
        \output_data_bus_0000_wide_signal  <= 32'b0;
        \output_data_bus_0001_wide_signal  <= 32'b0;
        \output_data_bus_0002_wide_signal  <= 32'b0;
        \output_data_bus_0003_wide_signal  <= 32'b0;
        \output_data_bus_0004_wide_signal  <= 32'b0;
        \output_data_bus_0005_wide_signal  <= 32'b0;
        \output_data_bus_0006_wide_signal  <= 32'b0;
        \output_data_bus_0007_wide_signal  <= 32'b0;
        \output_data_bus_0008_wide_signal  <= 32'b0;
        \output_data_bus_0009_wide_signal  <= 32'b0;
        \output_data_bus_0010_wide_signal  <= 32'b0;
        \output_data_bus_0011_wide_signal  <= 32'b0;
        \output_data_bus_0012_wide_signal  <= 32'b0;
        \output_data_bus_0013_wide_signal  <= 32'b0;
        \output_data_bus_0014_wide_signal  <= 32'b0;
        \output_data_bus_0015_wide_signal  <= 32'b0;
        \output_data_bus_0016_wide_signal  <= 32'b0;
        \output_data_bus_0017_wide_signal  <= 32'b0;
        \output_data_bus_0018_wide_signal  <= 32'b0;
        \output_data_bus_0019_wide_signal  <= 32'b0;
        \output_data_bus_0020_wide_signal  <= 32'b0;
        \output_data_bus_0021_wide_signal  <= 32'b0;
        \output_data_bus_0022_wide_signal  <= 32'b0;
        \output_data_bus_0023_wide_signal  <= 32'b0;
        \output_data_bus_0024_wide_signal  <= 32'b0;
        \output_data_bus_0025_wide_signal  <= 32'b0;
        \output_data_bus_0026_wide_signal  <= 32'b0;
        \output_data_bus_0027_wide_signal  <= 32'b0;
        \output_data_bus_0028_wide_signal  <= 32'b0;
        \output_data_bus_0029_wide_signal  <= 32'b0;
        \output_data_bus_0030_wide_signal  <= 32'b0;
        \output_data_bus_0031_wide_signal  <= 32'b0;
        \output_data_bus_0032_wide_signal  <= 32'b0;
        \output_data_bus_0033_wide_signal  <= 32'b0;
        \output_data_bus_0034_wide_signal  <= 32'b0;
        \output_data_bus_0035_wide_signal  <= 32'b0;
        \output_data_bus_0036_wide_signal  <= 32'b0;
        \output_data_bus_0037_wide_signal  <= 32'b0;
        \output_data_bus_0038_wide_signal  <= 32'b0;
        \output_data_bus_0039_wide_signal  <= 32'b0;
        \output_data_bus_0040_wide_signal  <= 32'b0;
        \output_data_bus_0041_wide_signal  <= 32'b0;
        \output_data_bus_0042_wide_signal  <= 32'b0;
        \output_data_bus_0043_wide_signal  <= 32'b0;
        \output_data_bus_0044_wide_signal  <= 32'b0;
        \output_data_bus_0045_wide_signal  <= 32'b0;
        \output_data_bus_0046_wide_signal  <= 32'b0;
        \output_data_bus_0047_wide_signal  <= 32'b0;
        \output_data_bus_0048_wide_signal  <= 32'b0;
        \output_data_bus_0049_wide_signal  <= 32'b0;
    end else begin
        \output_data_bus_0000_wide_signal  <= \input_data_bus_0000_wide_signal  + 32'd1;
        \output_data_bus_0001_wide_signal  <= \input_data_bus_0001_wide_signal  + 32'd1;
        \output_data_bus_0002_wide_signal  <= \input_data_bus_0002_wide_signal  + 32'd1;
        \output_data_bus_0003_wide_signal  <= \input_data_bus_0003_wide_signal  + 32'd1;
        \output_data_bus_0004_wide_signal  <= \input_data_bus_0004_wide_signal  + 32'd1;
        \output_data_bus_0005_wide_signal  <= \input_data_bus_0005_wide_signal  + 32'd1;
        \output_data_bus_0006_wide_signal  <= \input_data_bus_0006_wide_signal  + 32'd1;
        \output_data_bus_0007_wide_signal  <= \input_data_bus_0007_wide_signal  + 32'd1;
        \output_data_bus_0008_wide_signal  <= \input_data_bus_0008_wide_signal  + 32'd1;
        \output_data_bus_0009_wide_signal  <= \input_data_bus_0009_wide_signal  + 32'd1;
        \output_data_bus_0010_wide_signal  <= \input_data_bus_0010_wide_signal  + 32'd1;
        \output_data_bus_0011_wide_signal  <= \input_data_bus_0011_wide_signal  + 32'd1;
        \output_data_bus_0012_wide_signal  <= \input_data_bus_0012_wide_signal  + 32'd1;
        \output_data_bus_0013_wide_signal  <= \input_data_bus_0013_wide_signal  + 32'd1;
        \output_data_bus_0014_wide_signal  <= \input_data_bus_0014_wide_signal  + 32'd1;
        \output_data_bus_0015_wide_signal  <= \input_data_bus_0015_wide_signal  + 32'd1;
        \output_data_bus_0016_wide_signal  <= \input_data_bus_0016_wide_signal  + 32'd1;
        \output_data_bus_0017_wide_signal  <= \input_data_bus_0017_wide_signal  + 32'd1;
        \output_data_bus_0018_wide_signal  <= \input_data_bus_0018_wide_signal  + 32'd1;
        \output_data_bus_0019_wide_signal  <= \input_data_bus_0019_wide_signal  + 32'd1;
        \output_data_bus_0020_wide_signal  <= \input_data_bus_0020_wide_signal  + 32'd1;
        \output_data_bus_0021_wide_signal  <= \input_data_bus_0021_wide_signal  + 32'd1;
        \output_data_bus_0022_wide_signal  <= \input_data_bus_0022_wide_signal  + 32'd1;
        \output_data_bus_0023_wide_signal  <= \input_data_bus_0023_wide_signal  + 32'd1;
        \output_data_bus_0024_wide_signal  <= \input_data_bus_0024_wide_signal  + 32'd1;
        \output_data_bus_0025_wide_signal  <= \input_data_bus_0025_wide_signal  + 32'd1;
        \output_data_bus_0026_wide_signal  <= \input_data_bus_0026_wide_signal  + 32'd1;
        \output_data_bus_0027_wide_signal  <= \input_data_bus_0027_wide_signal  + 32'd1;
        \output_data_bus_0028_wide_signal  <= \input_data_bus_0028_wide_signal  + 32'd1;
        \output_data_bus_0029_wide_signal  <= \input_data_bus_0029_wide_signal  + 32'd1;
        \output_data_bus_0030_wide_signal  <= \input_data_bus_0030_wide_signal  + 32'd1;
        \output_data_bus_0031_wide_signal  <= \input_data_bus_0031_wide_signal  + 32'd1;
        \output_data_bus_0032_wide_signal  <= \input_data_bus_0032_wide_signal  + 32'd1;
        \output_data_bus_0033_wide_signal  <= \input_data_bus_0033_wide_signal  + 32'd1;
        \output_data_bus_0034_wide_signal  <= \input_data_bus_0034_wide_signal  + 32'd1;
        \output_data_bus_0035_wide_signal  <= \input_data_bus_0035_wide_signal  + 32'd1;
        \output_data_bus_0036_wide_signal  <= \input_data_bus_0036_wide_signal  + 32'd1;
        \output_data_bus_0037_wide_signal  <= \input_data_bus_0037_wide_signal  + 32'd1;
        \output_data_bus_0038_wide_signal  <= \input_data_bus_0038_wide_signal  + 32'd1;
        \output_data_bus_0039_wide_signal  <= \input_data_bus_0039_wide_signal  + 32'd1;
        \output_data_bus_0040_wide_signal  <= \input_data_bus_0040_wide_signal  + 32'd1;
        \output_data_bus_0041_wide_signal  <= \input_data_bus_0041_wide_signal  + 32'd1;
        \output_data_bus_0042_wide_signal  <= \input_data_bus_0042_wide_signal  + 32'd1;
        \output_data_bus_0043_wide_signal  <= \input_data_bus_0043_wide_signal  + 32'd1;
        \output_data_bus_0044_wide_signal  <= \input_data_bus_0044_wide_signal  + 32'd1;
        \output_data_bus_0045_wide_signal  <= \input_data_bus_0045_wide_signal  + 32'd1;
        \output_data_bus_0046_wide_signal  <= \input_data_bus_0046_wide_signal  + 32'd1;
        \output_data_bus_0047_wide_signal  <= \input_data_bus_0047_wide_signal  + 32'd1;
        \output_data_bus_0048_wide_signal  <= \input_data_bus_0048_wide_signal  + 32'd1;
        \output_data_bus_0049_wide_signal  <= \input_data_bus_0049_wide_signal  + 32'd1;
    end
end

endmodule
